* NGSPICE file created from MIPSpipeline.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

.subckt MIPSpipeline VGND VPWR clk current_pc[0] current_pc[10] current_pc[11] current_pc[12]
+ current_pc[13] current_pc[14] current_pc[15] current_pc[16] current_pc[17] current_pc[18]
+ current_pc[19] current_pc[1] current_pc[20] current_pc[21] current_pc[22] current_pc[23]
+ current_pc[24] current_pc[25] current_pc[26] current_pc[27] current_pc[28] current_pc[29]
+ current_pc[2] current_pc[30] current_pc[31] current_pc[3] current_pc[4] current_pc[5]
+ current_pc[6] current_pc[7] current_pc[8] current_pc[9] reset
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_131_ net40 _060_ VGND VGND VPWR VPWR PC4\[30\] sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_4_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_114_ net14 net15 _050_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__and3_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput7 net7 VGND VGND VPWR VPWR current_pc[15] sky130_fd_sc_hd__buf_2
Xoutput20 net20 VGND VGND VPWR VPWR current_pc[28] sky130_fd_sc_hd__buf_2
Xoutput31 net31 VGND VGND VPWR VPWR current_pc[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_130_ net21 net23 _055_ _058_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_113_ net14 _050_ net59 VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold20 net10 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR current_pc[29] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput8 net8 VGND VGND VPWR VPWR current_pc[16] sky130_fd_sc_hd__buf_2
Xoutput10 net10 VGND VGND VPWR VPWR current_pc[18] sky130_fd_sc_hd__buf_2
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_189_ clknet_2_1__leaf_clk PC4\[29\] _027_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_112_ net55 _050_ VGND VGND VPWR VPWR PC4\[22\] sky130_fd_sc_hd__xor2_1
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 net16 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net11 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput22 net22 VGND VGND VPWR VPWR current_pc[2] sky130_fd_sc_hd__buf_2
Xoutput9 net9 VGND VGND VPWR VPWR current_pc[17] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR current_pc[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_188_ clknet_2_1__leaf_clk PC4\[28\] _026_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_1
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_111_ net51 _048_ _050_ VGND VGND VPWR VPWR PC4\[21\] sky130_fd_sc_hd__o21ba_1
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold22 net15 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 net28 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput23 net23 VGND VGND VPWR VPWR current_pc[30] sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR current_pc[20] sky130_fd_sc_hd__buf_2
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_187_ clknet_2_1__leaf_clk PC4\[27\] _025_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_8
X_110_ _044_ _049_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__and2_1
Xhold12 net26 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 net21 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput24 net24 VGND VGND VPWR VPWR current_pc[31] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput13 net13 VGND VGND VPWR VPWR current_pc[21] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_186_ clknet_2_1__leaf_clk PC4\[26\] _024_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload1 clknet_2_1__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_8
X_169_ clknet_2_2__leaf_clk PC4\[9\] _007_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfrtp_1
Xhold13 net2 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 net19 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput14 net14 VGND VGND VPWR VPWR current_pc[22] sky130_fd_sc_hd__buf_2
Xoutput25 net25 VGND VGND VPWR VPWR current_pc[3] sky130_fd_sc_hd__buf_2
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_185_ clknet_2_3__leaf_clk PC4\[25\] _023_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload2 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_099_ net6 net7 net8 net9 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__and4_1
X_168_ clknet_2_2__leaf_clk PC4\[8\] _006_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfrtp_1
Xhold25 net12 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 net13 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR current_pc[23] sky130_fd_sc_hd__buf_2
Xoutput26 net26 VGND VGND VPWR VPWR current_pc[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_184_ clknet_2_3__leaf_clk PC4\[24\] _022_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_098_ net45 _041_ VGND VGND VPWR VPWR PC4\[16\] sky130_fd_sc_hd__xor2_1
X_167_ clknet_2_2__leaf_clk PC4\[7\] _005_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfrtp_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold15 net9 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput27 net27 VGND VGND VPWR VPWR current_pc[5] sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VPWR VPWR current_pc[24] sky130_fd_sc_hd__buf_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ clknet_2_3__leaf_clk PC4\[23\] _021_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_3_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_097_ net8 _041_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and2_1
X_166_ clknet_2_2__leaf_clk PC4\[6\] _004_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_19_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 net6 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_149_ net34 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__inv_2
Xoutput17 net17 VGND VGND VPWR VPWR current_pc[25] sky130_fd_sc_hd__buf_2
Xoutput28 net28 VGND VGND VPWR VPWR current_pc[6] sky130_fd_sc_hd__buf_2
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ clknet_2_3__leaf_clk PC4\[22\] _020_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_096_ net44 _040_ VGND VGND VPWR VPWR PC4\[15\] sky130_fd_sc_hd__xnor2_1
X_165_ clknet_2_2__leaf_clk PC4\[5\] _003_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold17 net17 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_148_ net32 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__inv_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput18 net18 VGND VGND VPWR VPWR current_pc[26] sky130_fd_sc_hd__buf_2
X_079_ net46 _030_ VGND VGND VPWR VPWR PC4\[8\] sky130_fd_sc_hd__xnor2_1
Xoutput29 net29 VGND VGND VPWR VPWR current_pc[7] sky130_fd_sc_hd__buf_2
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_181_ clknet_2_3__leaf_clk PC4\[21\] _019_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
X_095_ net6 net7 _039_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__and3_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_164_ clknet_2_3__leaf_clk PC4\[4\] _002_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfrtp_1
Xhold18 net14 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_147_ net32 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__inv_2
X_078_ _030_ _031_ VGND VGND VPWR VPWR PC4\[7\] sky130_fd_sc_hd__and2_1
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput19 net19 VGND VGND VPWR VPWR current_pc[27] sky130_fd_sc_hd__buf_2
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout32 net35 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
X_180_ clknet_2_2__leaf_clk PC4\[20\] _018_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
X_094_ net53 _039_ VGND VGND VPWR VPWR PC4\[14\] sky130_fd_sc_hd__xor2_1
X_163_ clknet_2_3__leaf_clk PC4\[3\] _001_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfrtp_1
Xhold19 net18 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_146_ net32 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_077_ net28 _064_ net29 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a21o_1
X_129_ _059_ _060_ VGND VGND VPWR VPWR PC4\[29\] sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout33 net35 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_093_ net6 _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2_1
X_162_ clknet_2_2__leaf_clk PC4\[2\] _000_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfrtp_1
Xinput1 reset VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_145_ net32 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__inv_2
X_076_ net28 net29 _064_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nand3_1
X_128_ net21 _055_ _058_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__and3_1
XFILLER_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout34 net35 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_4
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_161_ net33 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
X_092_ net42 _037_ VGND VGND VPWR VPWR PC4\[13\] sky130_fd_sc_hd__xor2_1
X_144_ net32 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__inv_2
X_075_ net48 _064_ VGND VGND VPWR VPWR PC4\[6\] sky130_fd_sc_hd__xor2_1
X_127_ _055_ _058_ net60 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout35 net1 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
X_160_ net33 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
X_091_ _064_ _032_ _038_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_143_ net32 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__inv_2
X_074_ _064_ _065_ VGND VGND VPWR VPWR PC4\[5\] sky130_fd_sc_hd__and2b_1
XFILLER_7_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_126_ net39 _057_ VGND VGND VPWR VPWR PC4\[28\] sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_3_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ net10 net11 net12 net13 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__and4_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_090_ net2 net3 net4 net5 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__and4_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_142_ net32 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
X_073_ net22 net25 net26 net27 VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__a31o_1
X_125_ net18 net19 net20 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_108_ _047_ _048_ VGND VGND VPWR VPWR PC4\[20\] sky130_fd_sc_hd__nor2_1
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_141_ net32 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
X_072_ net22 net25 net26 net27 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__and4_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_124_ _056_ _057_ VGND VGND VPWR VPWR PC4\[27\] sky130_fd_sc_hd__nor2_1
XMIPSpipeline_36 VGND VGND VPWR VPWR MIPSpipeline_36/HI current_pc[0] sky130_fd_sc_hd__conb_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_107_ net12 _046_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__and2_1
XFILLER_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_071_ net49 _062_ VGND VGND VPWR VPWR PC4\[4\] sky130_fd_sc_hd__xnor2_1
X_140_ net32 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_123_ net18 net19 _055_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__and3_1
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XMIPSpipeline_37 VGND VGND VPWR VPWR MIPSpipeline_37/HI current_pc[1] sky130_fd_sc_hd__conb_1
X_106_ net62 _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_070_ _062_ _063_ VGND VGND VPWR VPWR PC4\[3\] sky130_fd_sc_hd__and2_1
X_122_ net18 _055_ net61 VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_105_ _045_ _046_ VGND VGND VPWR VPWR PC4\[19\] sky130_fd_sc_hd__nor2_1
XFILLER_8_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_121_ net56 _055_ VGND VGND VPWR VPWR PC4\[26\] sky130_fd_sc_hd__xor2_1
X_104_ net10 net11 _044_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__and3_1
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ _054_ _055_ VGND VGND VPWR VPWR PC4\[25\] sky130_fd_sc_hd__nor2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_103_ net10 _044_ net58 VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 net24 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_179_ clknet_2_3__leaf_clk PC4\[19\] _017_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_102_ net57 _044_ VGND VGND VPWR VPWR PC4\[18\] sky130_fd_sc_hd__xor2_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 net20 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_178_ clknet_2_3__leaf_clk PC4\[18\] _016_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
X_101_ net52 _042_ _044_ VGND VGND VPWR VPWR PC4\[17\] sky130_fd_sc_hd__o21ba_1
Xhold3 net23 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_177_ clknet_2_0__leaf_clk PC4\[17\] _015_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
X_100_ _064_ _032_ _038_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__and4_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 net22 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_176_ clknet_2_1__leaf_clk PC4\[16\] _014_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_159_ net33 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 net5 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_175_ clknet_2_0__leaf_clk PC4\[15\] _013_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_089_ net43 _035_ VGND VGND VPWR VPWR PC4\[12\] sky130_fd_sc_hd__xor2_1
X_158_ net33 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__inv_2
XFILLER_8_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 net4 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_191_ clknet_2_1__leaf_clk PC4\[31\] _029_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfrtp_1
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_174_ clknet_2_0__leaf_clk PC4\[14\] _012_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfrtp_1
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_088_ net4 _035_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__and2_1
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_157_ net33 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__inv_2
Xhold7 net7 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ clknet_2_1__leaf_clk PC4\[30\] _028_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfrtp_1
X_173_ clknet_2_0__leaf_clk PC4\[13\] _011_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfrtp_1
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ _035_ _036_ VGND VGND VPWR VPWR PC4\[11\] sky130_fd_sc_hd__and2b_1
X_156_ net33 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__inv_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold8 net8 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
X_139_ net32 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__inv_2
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_172_ clknet_2_0__leaf_clk PC4\[12\] _010_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfrtp_1
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ net2 _064_ _032_ net3 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__a31o_1
X_155_ net35 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__inv_2
Xhold9 net30 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
X_069_ net22 net25 VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__or2_1
X_138_ net34 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__inv_2
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_171_ clknet_2_0__leaf_clk PC4\[11\] _009_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfrtp_1
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_085_ net2 net3 _033_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__and3_1
X_154_ net35 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__inv_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_068_ net22 net25 VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nand2_1
X_137_ net34 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__inv_2
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ clknet_2_0__leaf_clk PC4\[10\] _008_ VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dfrtp_1
X_153_ net35 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__inv_2
X_084_ net50 _033_ VGND VGND VPWR VPWR PC4\[10\] sky130_fd_sc_hd__xor2_1
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_136_ net34 VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__inv_2
X_067_ net34 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_119_ net17 _044_ _049_ _053_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__and4_2
Xoutput2 net2 VGND VGND VPWR VPWR current_pc[10] sky130_fd_sc_hd__buf_2
X_152_ net35 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__inv_2
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_083_ _033_ _034_ VGND VGND VPWR VPWR PC4\[9\] sky130_fd_sc_hd__and2b_1
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_066_ net41 VGND VGND VPWR VPWR PC4\[2\] sky130_fd_sc_hd__inv_2
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_135_ net34 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__inv_2
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_118_ _050_ _053_ net54 VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_12_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput3 net3 VGND VGND VPWR VPWR current_pc[11] sky130_fd_sc_hd__buf_2
XFILLER_15_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_082_ net28 net29 net30 _064_ net31 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__a41o_1
X_151_ net34 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__inv_2
X_134_ net34 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__inv_2
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_117_ _050_ _053_ _052_ net47 VGND VGND VPWR VPWR PC4\[24\] sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_5_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput4 net4 VGND VGND VPWR VPWR current_pc[12] sky130_fd_sc_hd__buf_2
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_081_ _064_ _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__and2_1
X_150_ net34 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_133_ net34 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ net14 net15 net16 VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput5 net5 VGND VGND VPWR VPWR current_pc[13] sky130_fd_sc_hd__buf_2
X_080_ net28 net29 net30 net31 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__and4_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_132_ net38 _061_ VGND VGND VPWR VPWR PC4\[31\] sky130_fd_sc_hd__xor2_1
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_115_ _051_ _052_ VGND VGND VPWR VPWR PC4\[23\] sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_16_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput6 net6 VGND VGND VPWR VPWR current_pc[14] sky130_fd_sc_hd__buf_2
Xoutput30 net30 VGND VGND VPWR VPWR current_pc[8] sky130_fd_sc_hd__buf_2
.ends

