VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MIPSpipeline
  CLASS BLOCK ;
  FOREIGN MIPSpipeline ;
  ORIGIN 0.000 0.000 ;
  SIZE 67.035 BY 77.755 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 76.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 72.080 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 74.580 72.080 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.480 -0.020 72.080 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 11.120 -0.020 12.920 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.120 -0.020 22.920 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.120 -0.020 32.920 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.120 -0.020 42.920 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.120 -0.020 52.920 76.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 16.480 72.080 18.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 26.480 72.080 28.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 36.480 72.080 38.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 46.480 72.080 48.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 56.480 72.080 58.280 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 72.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 68.780 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 71.280 68.780 72.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.180 3.280 68.780 72.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.620 -0.020 9.420 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 17.620 -0.020 19.420 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.620 -0.020 29.420 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.620 -0.020 39.420 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.620 -0.020 49.420 76.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.620 -0.020 59.420 76.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 12.980 72.080 14.780 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 22.980 72.080 24.780 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 32.980 72.080 34.780 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 42.980 72.080 44.780 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 52.980 72.080 54.780 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 62.980 72.080 64.780 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END clk
  PIN current_pc[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 63.035 13.640 67.035 14.240 ;
    END
  END current_pc[0]
  PIN current_pc[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END current_pc[10]
  PIN current_pc[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END current_pc[11]
  PIN current_pc[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END current_pc[12]
  PIN current_pc[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END current_pc[13]
  PIN current_pc[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END current_pc[14]
  PIN current_pc[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END current_pc[15]
  PIN current_pc[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END current_pc[16]
  PIN current_pc[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END current_pc[17]
  PIN current_pc[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 37.440 67.035 38.040 ;
    END
  END current_pc[18]
  PIN current_pc[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 40.840 67.035 41.440 ;
    END
  END current_pc[19]
  PIN current_pc[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 63.035 64.640 67.035 65.240 ;
    END
  END current_pc[1]
  PIN current_pc[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 47.640 67.035 48.240 ;
    END
  END current_pc[20]
  PIN current_pc[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 54.440 67.035 55.040 ;
    END
  END current_pc[21]
  PIN current_pc[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 61.240 67.035 61.840 ;
    END
  END current_pc[22]
  PIN current_pc[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 57.840 67.035 58.440 ;
    END
  END current_pc[23]
  PIN current_pc[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 51.040 67.035 51.640 ;
    END
  END current_pc[24]
  PIN current_pc[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 44.240 67.035 44.840 ;
    END
  END current_pc[25]
  PIN current_pc[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 30.640 67.035 31.240 ;
    END
  END current_pc[26]
  PIN current_pc[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 34.040 67.035 34.640 ;
    END
  END current_pc[27]
  PIN current_pc[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 27.240 67.035 27.840 ;
    END
  END current_pc[28]
  PIN current_pc[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 20.440 67.035 21.040 ;
    END
  END current_pc[29]
  PIN current_pc[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 73.755 22.910 77.755 ;
    END
  END current_pc[2]
  PIN current_pc[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 17.040 67.035 17.640 ;
    END
  END current_pc[30]
  PIN current_pc[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END current_pc[31]
  PIN current_pc[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 73.755 26.130 77.755 ;
    END
  END current_pc[3]
  PIN current_pc[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 73.755 32.570 77.755 ;
    END
  END current_pc[4]
  PIN current_pc[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 73.755 29.350 77.755 ;
    END
  END current_pc[5]
  PIN current_pc[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END current_pc[6]
  PIN current_pc[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END current_pc[7]
  PIN current_pc[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END current_pc[8]
  PIN current_pc[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END current_pc[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 63.035 23.840 67.035 24.440 ;
    END
  END reset
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 61.370 65.365 ;
      LAYER li1 ;
        RECT 5.520 10.795 61.180 65.365 ;
      LAYER met1 ;
        RECT 4.210 10.640 61.180 65.520 ;
      LAYER met2 ;
        RECT 4.230 73.475 22.350 74.530 ;
        RECT 23.190 73.475 25.570 74.530 ;
        RECT 26.410 73.475 28.790 74.530 ;
        RECT 29.630 73.475 32.010 74.530 ;
        RECT 32.850 73.475 61.080 74.530 ;
        RECT 4.230 4.280 61.080 73.475 ;
        RECT 4.230 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 44.890 4.280 ;
        RECT 45.730 4.000 61.080 4.280 ;
      LAYER met3 ;
        RECT 3.990 64.240 62.635 65.445 ;
        RECT 3.990 62.240 63.035 64.240 ;
        RECT 3.990 60.840 62.635 62.240 ;
        RECT 3.990 58.840 63.035 60.840 ;
        RECT 4.400 57.440 62.635 58.840 ;
        RECT 3.990 55.440 63.035 57.440 ;
        RECT 3.990 54.040 62.635 55.440 ;
        RECT 3.990 52.040 63.035 54.040 ;
        RECT 3.990 50.640 62.635 52.040 ;
        RECT 3.990 48.640 63.035 50.640 ;
        RECT 4.400 47.240 62.635 48.640 ;
        RECT 3.990 45.240 63.035 47.240 ;
        RECT 4.400 43.840 62.635 45.240 ;
        RECT 3.990 41.840 63.035 43.840 ;
        RECT 4.400 40.440 62.635 41.840 ;
        RECT 3.990 38.440 63.035 40.440 ;
        RECT 4.400 37.040 62.635 38.440 ;
        RECT 3.990 35.040 63.035 37.040 ;
        RECT 3.990 33.640 62.635 35.040 ;
        RECT 3.990 31.640 63.035 33.640 ;
        RECT 4.400 30.240 62.635 31.640 ;
        RECT 3.990 28.240 63.035 30.240 ;
        RECT 4.400 26.840 62.635 28.240 ;
        RECT 3.990 24.840 63.035 26.840 ;
        RECT 3.990 23.440 62.635 24.840 ;
        RECT 3.990 21.440 63.035 23.440 ;
        RECT 3.990 20.040 62.635 21.440 ;
        RECT 3.990 18.040 63.035 20.040 ;
        RECT 3.990 16.640 62.635 18.040 ;
        RECT 3.990 14.640 63.035 16.640 ;
        RECT 3.990 13.240 62.635 14.640 ;
        RECT 3.990 10.715 63.035 13.240 ;
  END
END MIPSpipeline
END LIBRARY

