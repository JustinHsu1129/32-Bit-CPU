module MIPSpipeline (clk,
    reset,
    current_pc);
 input clk;
 input reset;
 output [31:0] current_pc;

 wire \PC4[10] ;
 wire \PC4[11] ;
 wire \PC4[12] ;
 wire \PC4[13] ;
 wire \PC4[14] ;
 wire \PC4[15] ;
 wire \PC4[16] ;
 wire \PC4[17] ;
 wire \PC4[18] ;
 wire \PC4[19] ;
 wire \PC4[20] ;
 wire \PC4[21] ;
 wire \PC4[22] ;
 wire \PC4[23] ;
 wire \PC4[24] ;
 wire \PC4[25] ;
 wire \PC4[26] ;
 wire \PC4[27] ;
 wire \PC4[28] ;
 wire \PC4[29] ;
 wire \PC4[2] ;
 wire \PC4[30] ;
 wire \PC4[31] ;
 wire \PC4[3] ;
 wire \PC4[4] ;
 wire \PC4[5] ;
 wire \PC4[6] ;
 wire \PC4[7] ;
 wire \PC4[8] ;
 wire \PC4[9] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire net37;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;

 sky130_fd_sc_hd__inv_2 _066_ (.A(net41),
    .Y(\PC4[2] ));
 sky130_fd_sc_hd__inv_2 _067_ (.A(net34),
    .Y(_000_));
 sky130_fd_sc_hd__nand2_1 _068_ (.A(net22),
    .B(net25),
    .Y(_062_));
 sky130_fd_sc_hd__or2_1 _069_ (.A(net22),
    .B(net25),
    .X(_063_));
 sky130_fd_sc_hd__and2_1 _070_ (.A(_062_),
    .B(_063_),
    .X(\PC4[3] ));
 sky130_fd_sc_hd__xnor2_1 _071_ (.A(net49),
    .B(_062_),
    .Y(\PC4[4] ));
 sky130_fd_sc_hd__and4_2 _072_ (.A(net22),
    .B(net25),
    .C(net26),
    .D(net27),
    .X(_064_));
 sky130_fd_sc_hd__a31o_1 _073_ (.A1(net22),
    .A2(net25),
    .A3(net26),
    .B1(net27),
    .X(_065_));
 sky130_fd_sc_hd__and2b_1 _074_ (.A_N(_064_),
    .B(_065_),
    .X(\PC4[5] ));
 sky130_fd_sc_hd__xor2_1 _075_ (.A(net48),
    .B(_064_),
    .X(\PC4[6] ));
 sky130_fd_sc_hd__nand3_1 _076_ (.A(net28),
    .B(net29),
    .C(_064_),
    .Y(_030_));
 sky130_fd_sc_hd__a21o_1 _077_ (.A1(net28),
    .A2(_064_),
    .B1(net29),
    .X(_031_));
 sky130_fd_sc_hd__and2_1 _078_ (.A(_030_),
    .B(_031_),
    .X(\PC4[7] ));
 sky130_fd_sc_hd__xnor2_1 _079_ (.A(net46),
    .B(_030_),
    .Y(\PC4[8] ));
 sky130_fd_sc_hd__and4_1 _080_ (.A(net28),
    .B(net29),
    .C(net30),
    .D(net31),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _081_ (.A(_064_),
    .B(_032_),
    .X(_033_));
 sky130_fd_sc_hd__a41o_1 _082_ (.A1(net28),
    .A2(net29),
    .A3(net30),
    .A4(_064_),
    .B1(net31),
    .X(_034_));
 sky130_fd_sc_hd__and2b_1 _083_ (.A_N(_033_),
    .B(_034_),
    .X(\PC4[9] ));
 sky130_fd_sc_hd__xor2_1 _084_ (.A(net50),
    .B(_033_),
    .X(\PC4[10] ));
 sky130_fd_sc_hd__and3_1 _085_ (.A(net2),
    .B(net3),
    .C(_033_),
    .X(_035_));
 sky130_fd_sc_hd__a31o_1 _086_ (.A1(net2),
    .A2(_064_),
    .A3(_032_),
    .B1(net3),
    .X(_036_));
 sky130_fd_sc_hd__and2b_1 _087_ (.A_N(_035_),
    .B(_036_),
    .X(\PC4[11] ));
 sky130_fd_sc_hd__and2_1 _088_ (.A(net4),
    .B(_035_),
    .X(_037_));
 sky130_fd_sc_hd__xor2_1 _089_ (.A(net43),
    .B(_035_),
    .X(\PC4[12] ));
 sky130_fd_sc_hd__and4_1 _090_ (.A(net2),
    .B(net3),
    .C(net4),
    .D(net5),
    .X(_038_));
 sky130_fd_sc_hd__and3_1 _091_ (.A(_064_),
    .B(_032_),
    .C(_038_),
    .X(_039_));
 sky130_fd_sc_hd__xor2_1 _092_ (.A(net42),
    .B(_037_),
    .X(\PC4[13] ));
 sky130_fd_sc_hd__nand2_1 _093_ (.A(net6),
    .B(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__xor2_1 _094_ (.A(net53),
    .B(_039_),
    .X(\PC4[14] ));
 sky130_fd_sc_hd__and3_1 _095_ (.A(net6),
    .B(net7),
    .C(_039_),
    .X(_041_));
 sky130_fd_sc_hd__xnor2_1 _096_ (.A(net44),
    .B(_040_),
    .Y(\PC4[15] ));
 sky130_fd_sc_hd__and2_1 _097_ (.A(net8),
    .B(_041_),
    .X(_042_));
 sky130_fd_sc_hd__xor2_1 _098_ (.A(net45),
    .B(_041_),
    .X(\PC4[16] ));
 sky130_fd_sc_hd__and4_1 _099_ (.A(net6),
    .B(net7),
    .C(net8),
    .D(net9),
    .X(_043_));
 sky130_fd_sc_hd__and4_1 _100_ (.A(_064_),
    .B(_032_),
    .C(_038_),
    .D(_043_),
    .X(_044_));
 sky130_fd_sc_hd__o21ba_1 _101_ (.A1(net52),
    .A2(_042_),
    .B1_N(_044_),
    .X(\PC4[17] ));
 sky130_fd_sc_hd__xor2_1 _102_ (.A(net57),
    .B(_044_),
    .X(\PC4[18] ));
 sky130_fd_sc_hd__a21oi_1 _103_ (.A1(net10),
    .A2(_044_),
    .B1(net58),
    .Y(_045_));
 sky130_fd_sc_hd__and3_1 _104_ (.A(net10),
    .B(net11),
    .C(_044_),
    .X(_046_));
 sky130_fd_sc_hd__nor2_1 _105_ (.A(_045_),
    .B(_046_),
    .Y(\PC4[19] ));
 sky130_fd_sc_hd__nor2_1 _106_ (.A(net62),
    .B(_046_),
    .Y(_047_));
 sky130_fd_sc_hd__and2_1 _107_ (.A(net12),
    .B(_046_),
    .X(_048_));
 sky130_fd_sc_hd__nor2_1 _108_ (.A(_047_),
    .B(_048_),
    .Y(\PC4[20] ));
 sky130_fd_sc_hd__and4_1 _109_ (.A(net10),
    .B(net11),
    .C(net12),
    .D(net13),
    .X(_049_));
 sky130_fd_sc_hd__and2_1 _110_ (.A(_044_),
    .B(_049_),
    .X(_050_));
 sky130_fd_sc_hd__o21ba_1 _111_ (.A1(net51),
    .A2(_048_),
    .B1_N(_050_),
    .X(\PC4[21] ));
 sky130_fd_sc_hd__xor2_1 _112_ (.A(net55),
    .B(_050_),
    .X(\PC4[22] ));
 sky130_fd_sc_hd__a21oi_1 _113_ (.A1(net14),
    .A2(_050_),
    .B1(net59),
    .Y(_051_));
 sky130_fd_sc_hd__and3_1 _114_ (.A(net14),
    .B(net15),
    .C(_050_),
    .X(_052_));
 sky130_fd_sc_hd__nor2_1 _115_ (.A(_051_),
    .B(_052_),
    .Y(\PC4[23] ));
 sky130_fd_sc_hd__and3_1 _116_ (.A(net14),
    .B(net15),
    .C(net16),
    .X(_053_));
 sky130_fd_sc_hd__o2bb2a_1 _117_ (.A1_N(_050_),
    .A2_N(_053_),
    .B1(_052_),
    .B2(net47),
    .X(\PC4[24] ));
 sky130_fd_sc_hd__a21oi_1 _118_ (.A1(_050_),
    .A2(_053_),
    .B1(net54),
    .Y(_054_));
 sky130_fd_sc_hd__and4_2 _119_ (.A(net17),
    .B(_044_),
    .C(_049_),
    .D(_053_),
    .X(_055_));
 sky130_fd_sc_hd__nor2_1 _120_ (.A(_054_),
    .B(_055_),
    .Y(\PC4[25] ));
 sky130_fd_sc_hd__xor2_1 _121_ (.A(net56),
    .B(_055_),
    .X(\PC4[26] ));
 sky130_fd_sc_hd__a21oi_1 _122_ (.A1(net18),
    .A2(_055_),
    .B1(net61),
    .Y(_056_));
 sky130_fd_sc_hd__and3_1 _123_ (.A(net18),
    .B(net19),
    .C(_055_),
    .X(_057_));
 sky130_fd_sc_hd__nor2_1 _124_ (.A(_056_),
    .B(_057_),
    .Y(\PC4[27] ));
 sky130_fd_sc_hd__and3_1 _125_ (.A(net18),
    .B(net19),
    .C(net20),
    .X(_058_));
 sky130_fd_sc_hd__xor2_1 _126_ (.A(net39),
    .B(_057_),
    .X(\PC4[28] ));
 sky130_fd_sc_hd__a21oi_1 _127_ (.A1(_055_),
    .A2(_058_),
    .B1(net60),
    .Y(_059_));
 sky130_fd_sc_hd__and3_1 _128_ (.A(net21),
    .B(_055_),
    .C(_058_),
    .X(_060_));
 sky130_fd_sc_hd__nor2_1 _129_ (.A(_059_),
    .B(_060_),
    .Y(\PC4[29] ));
 sky130_fd_sc_hd__and4_1 _130_ (.A(net21),
    .B(net23),
    .C(_055_),
    .D(_058_),
    .X(_061_));
 sky130_fd_sc_hd__xor2_1 _131_ (.A(net40),
    .B(_060_),
    .X(\PC4[30] ));
 sky130_fd_sc_hd__xor2_1 _132_ (.A(net38),
    .B(_061_),
    .X(\PC4[31] ));
 sky130_fd_sc_hd__inv_2 _133_ (.A(net34),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _134_ (.A(net34),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _135_ (.A(net34),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _136_ (.A(net34),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _137_ (.A(net34),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _138_ (.A(net34),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _139_ (.A(net32),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _140_ (.A(net32),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _141_ (.A(net32),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _142_ (.A(net32),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _143_ (.A(net32),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _144_ (.A(net32),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _145_ (.A(net32),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _146_ (.A(net32),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _147_ (.A(net32),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _148_ (.A(net32),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _149_ (.A(net34),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _150_ (.A(net34),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _151_ (.A(net34),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _152_ (.A(net35),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _153_ (.A(net35),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _154_ (.A(net35),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _155_ (.A(net35),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _156_ (.A(net33),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _157_ (.A(net33),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _158_ (.A(net33),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _159_ (.A(net33),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _160_ (.A(net33),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _161_ (.A(net33),
    .Y(_029_));
 sky130_fd_sc_hd__dfrtp_1 _162_ (.CLK(clknet_2_2__leaf_clk),
    .D(\PC4[2] ),
    .RESET_B(_000_),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _163_ (.CLK(clknet_2_3__leaf_clk),
    .D(\PC4[3] ),
    .RESET_B(_001_),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _164_ (.CLK(clknet_2_3__leaf_clk),
    .D(\PC4[4] ),
    .RESET_B(_002_),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _165_ (.CLK(clknet_2_2__leaf_clk),
    .D(\PC4[5] ),
    .RESET_B(_003_),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_2 _166_ (.CLK(clknet_2_2__leaf_clk),
    .D(\PC4[6] ),
    .RESET_B(_004_),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _167_ (.CLK(clknet_2_2__leaf_clk),
    .D(\PC4[7] ),
    .RESET_B(_005_),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _168_ (.CLK(clknet_2_2__leaf_clk),
    .D(\PC4[8] ),
    .RESET_B(_006_),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _169_ (.CLK(clknet_2_2__leaf_clk),
    .D(\PC4[9] ),
    .RESET_B(_007_),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _170_ (.CLK(clknet_2_0__leaf_clk),
    .D(\PC4[10] ),
    .RESET_B(_008_),
    .Q(net2));
 sky130_fd_sc_hd__dfrtp_1 _171_ (.CLK(clknet_2_0__leaf_clk),
    .D(\PC4[11] ),
    .RESET_B(_009_),
    .Q(net3));
 sky130_fd_sc_hd__dfrtp_1 _172_ (.CLK(clknet_2_0__leaf_clk),
    .D(\PC4[12] ),
    .RESET_B(_010_),
    .Q(net4));
 sky130_fd_sc_hd__dfrtp_1 _173_ (.CLK(clknet_2_0__leaf_clk),
    .D(\PC4[13] ),
    .RESET_B(_011_),
    .Q(net5));
 sky130_fd_sc_hd__dfrtp_1 _174_ (.CLK(clknet_2_0__leaf_clk),
    .D(\PC4[14] ),
    .RESET_B(_012_),
    .Q(net6));
 sky130_fd_sc_hd__dfrtp_1 _175_ (.CLK(clknet_2_0__leaf_clk),
    .D(\PC4[15] ),
    .RESET_B(_013_),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_1 _176_ (.CLK(clknet_2_1__leaf_clk),
    .D(\PC4[16] ),
    .RESET_B(_014_),
    .Q(net8));
 sky130_fd_sc_hd__dfrtp_1 _177_ (.CLK(clknet_2_0__leaf_clk),
    .D(\PC4[17] ),
    .RESET_B(_015_),
    .Q(net9));
 sky130_fd_sc_hd__dfrtp_1 _178_ (.CLK(clknet_2_3__leaf_clk),
    .D(\PC4[18] ),
    .RESET_B(_016_),
    .Q(net10));
 sky130_fd_sc_hd__dfrtp_1 _179_ (.CLK(clknet_2_3__leaf_clk),
    .D(\PC4[19] ),
    .RESET_B(_017_),
    .Q(net11));
 sky130_fd_sc_hd__dfrtp_1 _180_ (.CLK(clknet_2_2__leaf_clk),
    .D(\PC4[20] ),
    .RESET_B(_018_),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_1 _181_ (.CLK(clknet_2_3__leaf_clk),
    .D(\PC4[21] ),
    .RESET_B(_019_),
    .Q(net13));
 sky130_fd_sc_hd__dfrtp_1 _182_ (.CLK(clknet_2_3__leaf_clk),
    .D(\PC4[22] ),
    .RESET_B(_020_),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_1 _183_ (.CLK(clknet_2_3__leaf_clk),
    .D(\PC4[23] ),
    .RESET_B(_021_),
    .Q(net15));
 sky130_fd_sc_hd__dfrtp_1 _184_ (.CLK(clknet_2_3__leaf_clk),
    .D(\PC4[24] ),
    .RESET_B(_022_),
    .Q(net16));
 sky130_fd_sc_hd__dfrtp_1 _185_ (.CLK(clknet_2_3__leaf_clk),
    .D(\PC4[25] ),
    .RESET_B(_023_),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_1 _186_ (.CLK(clknet_2_1__leaf_clk),
    .D(\PC4[26] ),
    .RESET_B(_024_),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_1 _187_ (.CLK(clknet_2_1__leaf_clk),
    .D(\PC4[27] ),
    .RESET_B(_025_),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 _188_ (.CLK(clknet_2_1__leaf_clk),
    .D(\PC4[28] ),
    .RESET_B(_026_),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _189_ (.CLK(clknet_2_1__leaf_clk),
    .D(\PC4[29] ),
    .RESET_B(_027_),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _190_ (.CLK(clknet_2_1__leaf_clk),
    .D(\PC4[30] ),
    .RESET_B(_028_),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _191_ (.CLK(clknet_2_1__leaf_clk),
    .D(\PC4[31] ),
    .RESET_B(_029_),
    .Q(net24));
 sky130_fd_sc_hd__conb_1 MIPSpipeline_37 (.LO(net37));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_83 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(reset),
    .X(net1));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(current_pc[10]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(current_pc[11]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(current_pc[12]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(current_pc[13]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(current_pc[14]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(current_pc[15]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(current_pc[16]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(current_pc[17]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(current_pc[18]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(current_pc[19]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(current_pc[20]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(current_pc[21]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(current_pc[22]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(current_pc[23]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(current_pc[24]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(current_pc[25]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(current_pc[26]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(current_pc[27]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(current_pc[28]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(current_pc[29]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(current_pc[2]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(current_pc[30]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(current_pc[31]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(current_pc[3]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(current_pc[4]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(current_pc[5]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(current_pc[6]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(current_pc[7]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(current_pc[8]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(current_pc[9]));
 sky130_fd_sc_hd__buf_4 fanout32 (.A(net35),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(net35),
    .X(net33));
 sky130_fd_sc_hd__buf_4 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(net1),
    .X(net35));
 sky130_fd_sc_hd__conb_1 MIPSpipeline_36 (.LO(net36));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload1 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net24),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net20),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net23),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net22),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net5),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net4),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net7),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net8),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net30),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net16),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net28),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net26),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net2),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net13),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net9),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net6),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net17),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net14),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net18),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net10),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net11),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net15),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net21),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net19),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net12),
    .X(net62));
 assign current_pc[0] = net36;
 assign current_pc[1] = net37;
endmodule
