magic
tech sky130A
magscale 1 2
timestamp 1757946788
<< viali >>
rect 4537 12937 4571 12971
rect 4997 12937 5031 12971
rect 6101 12937 6135 12971
rect 6745 12937 6779 12971
rect 9873 12869 9907 12903
rect 4721 12801 4755 12835
rect 4813 12801 4847 12835
rect 5365 12801 5399 12835
rect 5917 12801 5951 12835
rect 6561 12801 6595 12835
rect 9781 12801 9815 12835
rect 10057 12801 10091 12835
rect 10241 12801 10275 12835
rect 10333 12801 10367 12835
rect 11621 12801 11655 12835
rect 5457 12733 5491 12767
rect 10701 12733 10735 12767
rect 5733 12665 5767 12699
rect 9689 12665 9723 12699
rect 10057 12597 10091 12631
rect 10517 12597 10551 12631
rect 11345 12597 11379 12631
rect 11805 12597 11839 12631
rect 5457 12393 5491 12427
rect 5917 12393 5951 12427
rect 10057 12393 10091 12427
rect 9873 12325 9907 12359
rect 10333 12325 10367 12359
rect 5181 12257 5215 12291
rect 6561 12257 6595 12291
rect 10885 12257 10919 12291
rect 11161 12257 11195 12291
rect 3985 12189 4019 12223
rect 4445 12189 4479 12223
rect 4629 12189 4663 12223
rect 5365 12189 5399 12223
rect 5549 12189 5583 12223
rect 6837 12189 6871 12223
rect 7113 12189 7147 12223
rect 9413 12189 9447 12223
rect 10458 12189 10492 12223
rect 10977 12189 11011 12223
rect 11713 12189 11747 12223
rect 6653 12121 6687 12155
rect 10241 12121 10275 12155
rect 4077 12053 4111 12087
rect 4353 12053 4387 12087
rect 7021 12053 7055 12087
rect 7205 12053 7239 12087
rect 9505 12053 9539 12087
rect 10041 12053 10075 12087
rect 10517 12053 10551 12087
rect 3341 11781 3375 11815
rect 11345 11781 11379 11815
rect 5273 11713 5307 11747
rect 5365 11713 5399 11747
rect 5457 11713 5491 11747
rect 5733 11713 5767 11747
rect 5917 11713 5951 11747
rect 11069 11713 11103 11747
rect 11161 11713 11195 11747
rect 11621 11713 11655 11747
rect 3065 11645 3099 11679
rect 7849 11645 7883 11679
rect 8125 11645 8159 11679
rect 8493 11645 8527 11679
rect 8769 11645 8803 11679
rect 10241 11645 10275 11679
rect 10977 11645 11011 11679
rect 4813 11577 4847 11611
rect 5641 11577 5675 11611
rect 6377 11577 6411 11611
rect 10333 11577 10367 11611
rect 11345 11577 11379 11611
rect 5089 11509 5123 11543
rect 6101 11509 6135 11543
rect 11805 11509 11839 11543
rect 4629 11305 4663 11339
rect 5273 11305 5307 11339
rect 8953 11305 8987 11339
rect 11897 11305 11931 11339
rect 4353 11237 4387 11271
rect 3985 11169 4019 11203
rect 4445 11169 4479 11203
rect 4813 11169 4847 11203
rect 5089 11169 5123 11203
rect 6745 11169 6779 11203
rect 9229 11169 9263 11203
rect 10425 11169 10459 11203
rect 4905 11101 4939 11135
rect 4997 11101 5031 11135
rect 7021 11101 7055 11135
rect 7297 11101 7331 11135
rect 9321 11101 9355 11135
rect 10149 11101 10183 11135
rect 7205 11033 7239 11067
rect 5641 10761 5675 10795
rect 11345 10761 11379 10795
rect 11729 10761 11763 10795
rect 11897 10761 11931 10795
rect 11529 10693 11563 10727
rect 1685 10625 1719 10659
rect 3893 10625 3927 10659
rect 8493 10625 8527 10659
rect 9505 10625 9539 10659
rect 9597 10625 9631 10659
rect 4169 10557 4203 10591
rect 8677 10557 8711 10591
rect 9873 10557 9907 10591
rect 1501 10421 1535 10455
rect 8309 10421 8343 10455
rect 9413 10421 9447 10455
rect 11713 10421 11747 10455
rect 4905 10217 4939 10251
rect 11621 10217 11655 10251
rect 1501 10081 1535 10115
rect 1961 10081 1995 10115
rect 3157 10081 3191 10115
rect 1869 10013 1903 10047
rect 2605 10013 2639 10047
rect 3525 10013 3559 10047
rect 3985 10013 4019 10047
rect 4169 10013 4203 10047
rect 4813 10013 4847 10047
rect 7849 10013 7883 10047
rect 8033 10013 8067 10047
rect 8309 10013 8343 10047
rect 8585 10013 8619 10047
rect 8769 10013 8803 10047
rect 10977 10013 11011 10047
rect 11437 10013 11471 10047
rect 3801 9945 3835 9979
rect 8953 9945 8987 9979
rect 11069 9945 11103 9979
rect 11345 9945 11379 9979
rect 3433 9877 3467 9911
rect 7941 9877 7975 9911
rect 8125 9877 8159 9911
rect 10241 9877 10275 9911
rect 10793 9877 10827 9911
rect 11161 9877 11195 9911
rect 3249 9673 3283 9707
rect 1777 9605 1811 9639
rect 5549 9605 5583 9639
rect 9781 9605 9815 9639
rect 11713 9605 11747 9639
rect 7665 9537 7699 9571
rect 10425 9537 10459 9571
rect 11345 9537 11379 9571
rect 11529 9537 11563 9571
rect 11805 9537 11839 9571
rect 1501 9469 1535 9503
rect 7941 9469 7975 9503
rect 8217 9469 8251 9503
rect 9689 9469 9723 9503
rect 10793 9469 10827 9503
rect 11529 9401 11563 9435
rect 4077 9333 4111 9367
rect 7757 9333 7791 9367
rect 5549 9129 5583 9163
rect 6101 9129 6135 9163
rect 8769 9129 8803 9163
rect 10057 9129 10091 9163
rect 1501 9061 1535 9095
rect 1869 9061 1903 9095
rect 6561 9061 6595 9095
rect 3617 8993 3651 9027
rect 7021 8993 7055 9027
rect 7297 8993 7331 9027
rect 9505 8993 9539 9027
rect 10149 8993 10183 9027
rect 1685 8925 1719 8959
rect 3801 8925 3835 8959
rect 5365 8925 5399 8959
rect 5733 8925 5767 8959
rect 6009 8925 6043 8959
rect 6101 8925 6135 8959
rect 6653 8925 6687 8959
rect 9781 8925 9815 8959
rect 9873 8925 9907 8959
rect 3341 8857 3375 8891
rect 6193 8857 6227 8891
rect 6377 8857 6411 8891
rect 10425 8857 10459 8891
rect 4813 8789 4847 8823
rect 5917 8789 5951 8823
rect 8953 8789 8987 8823
rect 11897 8789 11931 8823
rect 2237 8585 2271 8619
rect 2421 8585 2455 8619
rect 5549 8585 5583 8619
rect 7941 8585 7975 8619
rect 9781 8585 9815 8619
rect 10609 8585 10643 8619
rect 11805 8585 11839 8619
rect 5733 8517 5767 8551
rect 9933 8517 9967 8551
rect 10149 8517 10183 8551
rect 10885 8517 10919 8551
rect 1685 8449 1719 8483
rect 2513 8449 2547 8483
rect 3249 8449 3283 8483
rect 3801 8449 3835 8483
rect 5825 8449 5859 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 7849 8449 7883 8483
rect 8125 8449 8159 8483
rect 8493 8449 8527 8483
rect 9229 8449 9263 8483
rect 10517 8449 10551 8483
rect 10701 8449 10735 8483
rect 11069 8449 11103 8483
rect 11621 8449 11655 8483
rect 2053 8381 2087 8415
rect 2145 8381 2179 8415
rect 3341 8381 3375 8415
rect 4077 8381 4111 8415
rect 9045 8381 9079 8415
rect 9505 8381 9539 8415
rect 1501 8313 1535 8347
rect 1869 8313 1903 8347
rect 3617 8313 3651 8347
rect 8125 8313 8159 8347
rect 11253 8313 11287 8347
rect 7573 8245 7607 8279
rect 9965 8245 9999 8279
rect 10333 8245 10367 8279
rect 6653 8041 6687 8075
rect 8953 8041 8987 8075
rect 9413 8041 9447 8075
rect 10793 8041 10827 8075
rect 11069 8041 11103 8075
rect 11805 8041 11839 8075
rect 2329 7973 2363 8007
rect 8769 7973 8803 8007
rect 7297 7905 7331 7939
rect 1685 7837 1719 7871
rect 5181 7837 5215 7871
rect 7021 7837 7055 7871
rect 8953 7837 8987 7871
rect 9137 7837 9171 7871
rect 9413 7837 9447 7871
rect 9597 7837 9631 7871
rect 9689 7837 9723 7871
rect 10701 7837 10735 7871
rect 11161 7837 11195 7871
rect 11253 7837 11287 7871
rect 11621 7837 11655 7871
rect 2513 7769 2547 7803
rect 2605 7769 2639 7803
rect 9781 7769 9815 7803
rect 1501 7701 1535 7735
rect 2697 7701 2731 7735
rect 2881 7701 2915 7735
rect 11437 7701 11471 7735
rect 3249 7497 3283 7531
rect 8769 7497 8803 7531
rect 3433 7429 3467 7463
rect 9689 7429 9723 7463
rect 1501 7361 1535 7395
rect 3525 7361 3559 7395
rect 7021 7361 7055 7395
rect 9413 7361 9447 7395
rect 9597 7361 9631 7395
rect 10425 7361 10459 7395
rect 11529 7361 11563 7395
rect 1777 7293 1811 7327
rect 7297 7293 7331 7327
rect 10793 7293 10827 7327
rect 8861 7225 8895 7259
rect 10517 7157 10551 7191
rect 11345 7157 11379 7191
rect 11713 7157 11747 7191
rect 1777 6953 1811 6987
rect 7113 6953 7147 6987
rect 1869 6885 1903 6919
rect 7389 6817 7423 6851
rect 8953 6817 8987 6851
rect 9413 6817 9447 6851
rect 7481 6749 7515 6783
rect 9321 6749 9355 6783
rect 9965 6749 9999 6783
rect 2237 6681 2271 6715
rect 10241 6681 10275 6715
rect 11713 6613 11747 6647
rect 8861 6409 8895 6443
rect 1961 6341 1995 6375
rect 2161 6341 2195 6375
rect 3249 6341 3283 6375
rect 4905 6341 4939 6375
rect 5105 6341 5139 6375
rect 1685 6273 1719 6307
rect 3433 6273 3467 6307
rect 3525 6273 3559 6307
rect 3893 6273 3927 6307
rect 3985 6273 4019 6307
rect 9597 6273 9631 6307
rect 11529 6273 11563 6307
rect 2697 6205 2731 6239
rect 9413 6205 9447 6239
rect 3065 6137 3099 6171
rect 1501 6069 1535 6103
rect 2145 6069 2179 6103
rect 2329 6069 2363 6103
rect 3157 6069 3191 6103
rect 3801 6069 3835 6103
rect 4077 6069 4111 6103
rect 5089 6069 5123 6103
rect 5273 6069 5307 6103
rect 9860 6069 9894 6103
rect 11345 6069 11379 6103
rect 11713 6069 11747 6103
rect 3617 5865 3651 5899
rect 9965 5865 9999 5899
rect 11621 5797 11655 5831
rect 5273 5729 5307 5763
rect 10425 5729 10459 5763
rect 11437 5729 11471 5763
rect 1685 5661 1719 5695
rect 1869 5661 1903 5695
rect 5549 5661 5583 5695
rect 5641 5661 5675 5695
rect 8033 5661 8067 5695
rect 8401 5661 8435 5695
rect 8769 5661 8803 5695
rect 10333 5661 10367 5695
rect 10885 5661 10919 5695
rect 11897 5661 11931 5695
rect 2145 5593 2179 5627
rect 5917 5593 5951 5627
rect 8953 5593 8987 5627
rect 11621 5593 11655 5627
rect 1501 5525 1535 5559
rect 3801 5525 3835 5559
rect 7389 5525 7423 5559
rect 7481 5525 7515 5559
rect 8309 5525 8343 5559
rect 8677 5525 8711 5559
rect 11805 5525 11839 5559
rect 3893 5321 3927 5355
rect 3985 5321 4019 5355
rect 4261 5321 4295 5355
rect 5549 5321 5583 5355
rect 6377 5321 6411 5355
rect 9689 5321 9723 5355
rect 9873 5321 9907 5355
rect 10425 5321 10459 5355
rect 11687 5321 11721 5355
rect 5457 5253 5491 5287
rect 5825 5253 5859 5287
rect 10777 5253 10811 5287
rect 10977 5253 11011 5287
rect 11897 5253 11931 5287
rect 1685 5185 1719 5219
rect 2697 5185 2731 5219
rect 3249 5185 3283 5219
rect 3709 5185 3743 5219
rect 4077 5185 4111 5219
rect 5273 5185 5307 5219
rect 5641 5185 5675 5219
rect 6561 5185 6595 5219
rect 6837 5185 6871 5219
rect 7021 5185 7055 5219
rect 7941 5185 7975 5219
rect 9781 5185 9815 5219
rect 9965 5185 9999 5219
rect 10057 5185 10091 5219
rect 10241 5185 10275 5219
rect 10333 5185 10367 5219
rect 11345 5185 11379 5219
rect 1777 5117 1811 5151
rect 2053 5117 2087 5151
rect 8217 5117 8251 5151
rect 10609 5049 10643 5083
rect 10241 4981 10275 5015
rect 10793 4981 10827 5015
rect 11161 4981 11195 5015
rect 11529 4981 11563 5015
rect 11713 4981 11747 5015
rect 3065 4777 3099 4811
rect 10241 4777 10275 4811
rect 10977 4777 11011 4811
rect 11805 4777 11839 4811
rect 11437 4709 11471 4743
rect 3249 4641 3283 4675
rect 3433 4641 3467 4675
rect 3525 4641 3559 4675
rect 6193 4641 6227 4675
rect 6653 4641 6687 4675
rect 6745 4641 6779 4675
rect 8493 4641 8527 4675
rect 3341 4573 3375 4607
rect 3985 4573 4019 4607
rect 4077 4573 4111 4607
rect 6285 4573 6319 4607
rect 11253 4573 11287 4607
rect 11621 4573 11655 4607
rect 4261 4505 4295 4539
rect 6009 4505 6043 4539
rect 7021 4505 7055 4539
rect 8953 4505 8987 4539
rect 11161 4505 11195 4539
rect 3801 4437 3835 4471
rect 10793 4437 10827 4471
rect 10961 4437 10995 4471
rect 5641 4233 5675 4267
rect 5825 4233 5859 4267
rect 9413 4233 9447 4267
rect 9505 4233 9539 4267
rect 9597 4233 9631 4267
rect 6009 4165 6043 4199
rect 9137 4165 9171 4199
rect 10609 4165 10643 4199
rect 2329 4097 2363 4131
rect 3525 4097 3559 4131
rect 4261 4097 4295 4131
rect 5549 4097 5583 4131
rect 5917 4097 5951 4131
rect 7389 4097 7423 4131
rect 8033 4097 8067 4131
rect 8585 4097 8619 4131
rect 8861 4097 8895 4131
rect 8953 4097 8987 4131
rect 9781 4097 9815 4131
rect 11161 4097 11195 4131
rect 11621 4097 11655 4131
rect 2421 4029 2455 4063
rect 3433 4029 3467 4063
rect 4077 4029 4111 4063
rect 6929 4029 6963 4063
rect 8401 4029 8435 4063
rect 9064 4029 9098 4063
rect 10425 4029 10459 4063
rect 6193 3961 6227 3995
rect 11805 3961 11839 3995
rect 2697 3893 2731 3927
rect 2789 3893 2823 3927
rect 5457 3893 5491 3927
rect 6377 3893 6411 3927
rect 9229 3893 9263 3927
rect 9873 3893 9907 3927
rect 7849 3689 7883 3723
rect 8033 3689 8067 3723
rect 8493 3689 8527 3723
rect 11437 3689 11471 3723
rect 1869 3553 1903 3587
rect 4169 3553 4203 3587
rect 6009 3553 6043 3587
rect 7757 3553 7791 3587
rect 9321 3553 9355 3587
rect 9597 3553 9631 3587
rect 9689 3553 9723 3587
rect 3985 3485 4019 3519
rect 8585 3485 8619 3519
rect 9229 3485 9263 3519
rect 11621 3485 11655 3519
rect 2145 3417 2179 3451
rect 3893 3417 3927 3451
rect 4445 3417 4479 3451
rect 6285 3417 6319 3451
rect 8217 3417 8251 3451
rect 9965 3417 9999 3451
rect 3617 3349 3651 3383
rect 5917 3349 5951 3383
rect 8007 3349 8041 3383
rect 11805 3349 11839 3383
rect 4629 3145 4663 3179
rect 6745 3145 6779 3179
rect 11529 3145 11563 3179
rect 3157 3077 3191 3111
rect 2329 3009 2363 3043
rect 2881 3009 2915 3043
rect 5273 3009 5307 3043
rect 5733 3009 5767 3043
rect 6561 3009 6595 3043
rect 7389 3009 7423 3043
rect 7665 3009 7699 3043
rect 9597 3009 9631 3043
rect 11713 3009 11747 3043
rect 1961 2941 1995 2975
rect 2421 2941 2455 2975
rect 4905 2941 4939 2975
rect 5365 2941 5399 2975
rect 5825 2941 5859 2975
rect 6377 2941 6411 2975
rect 6837 2941 6871 2975
rect 7941 2941 7975 2975
rect 9873 2941 9907 2975
rect 11345 2873 11379 2907
rect 6009 2805 6043 2839
rect 9413 2805 9447 2839
rect 4445 2601 4479 2635
rect 7021 2601 7055 2635
rect 7665 2601 7699 2635
rect 8217 2601 8251 2635
rect 9045 2601 9079 2635
rect 10977 2601 11011 2635
rect 11253 2601 11287 2635
rect 11897 2601 11931 2635
rect 8677 2465 8711 2499
rect 9965 2465 9999 2499
rect 3617 2397 3651 2431
rect 4261 2397 4295 2431
rect 4537 2397 4571 2431
rect 6193 2397 6227 2431
rect 6837 2397 6871 2431
rect 6929 2397 6963 2431
rect 7113 2397 7147 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 8125 2397 8159 2431
rect 8585 2397 8619 2431
rect 9137 2397 9171 2431
rect 10149 2397 10183 2431
rect 11069 2397 11103 2431
rect 11161 2397 11195 2431
rect 9413 2329 9447 2363
rect 3433 2261 3467 2295
rect 4077 2261 4111 2295
rect 6009 2261 6043 2295
rect 6653 2261 6687 2295
rect 7297 2261 7331 2295
rect 7941 2261 7975 2295
rect 10333 2261 10367 2295
<< metal1 >>
rect 1104 13082 12236 13104
rect 1104 13030 2250 13082
rect 2302 13030 2314 13082
rect 2366 13030 2378 13082
rect 2430 13030 2442 13082
rect 2494 13030 2506 13082
rect 2558 13030 4250 13082
rect 4302 13030 4314 13082
rect 4366 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 6250 13082
rect 6302 13030 6314 13082
rect 6366 13030 6378 13082
rect 6430 13030 6442 13082
rect 6494 13030 6506 13082
rect 6558 13030 8250 13082
rect 8302 13030 8314 13082
rect 8366 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 10250 13082
rect 10302 13030 10314 13082
rect 10366 13030 10378 13082
rect 10430 13030 10442 13082
rect 10494 13030 10506 13082
rect 10558 13030 12236 13082
rect 1104 13008 12236 13030
rect 4525 12971 4583 12977
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 4614 12968 4620 12980
rect 4571 12940 4620 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 4982 12928 4988 12980
rect 5040 12928 5046 12980
rect 6086 12928 6092 12980
rect 6144 12928 6150 12980
rect 6730 12928 6736 12980
rect 6788 12928 6794 12980
rect 9861 12903 9919 12909
rect 9861 12869 9873 12903
rect 9907 12900 9919 12903
rect 11054 12900 11060 12912
rect 9907 12872 11060 12900
rect 9907 12869 9919 12872
rect 9861 12863 9919 12869
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12832 4859 12835
rect 5258 12832 5264 12844
rect 4847 12804 5264 12832
rect 4847 12801 4859 12804
rect 4801 12795 4859 12801
rect 4724 12764 4752 12795
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5810 12832 5816 12844
rect 5399 12804 5816 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 5905 12835 5963 12841
rect 5905 12801 5917 12835
rect 5951 12832 5963 12835
rect 5994 12832 6000 12844
rect 5951 12804 6000 12832
rect 5951 12801 5963 12804
rect 5905 12795 5963 12801
rect 5994 12792 6000 12804
rect 6052 12792 6058 12844
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12832 6607 12835
rect 6638 12832 6644 12844
rect 6595 12804 6644 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12832 9827 12835
rect 9950 12832 9956 12844
rect 9815 12804 9956 12832
rect 9815 12801 9827 12804
rect 9769 12795 9827 12801
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 10042 12792 10048 12844
rect 10100 12792 10106 12844
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 5166 12764 5172 12776
rect 4724 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5442 12724 5448 12776
rect 5500 12724 5506 12776
rect 10244 12764 10272 12795
rect 10318 12792 10324 12844
rect 10376 12792 10382 12844
rect 11238 12832 11244 12844
rect 10612 12804 11244 12832
rect 10612 12764 10640 12804
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11609 12835 11667 12841
rect 11609 12801 11621 12835
rect 11655 12832 11667 12835
rect 12066 12832 12072 12844
rect 11655 12804 12072 12832
rect 11655 12801 11667 12804
rect 11609 12795 11667 12801
rect 10244 12736 10640 12764
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 11624 12764 11652 12795
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 10735 12736 11652 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 5721 12699 5779 12705
rect 5721 12665 5733 12699
rect 5767 12696 5779 12699
rect 7374 12696 7380 12708
rect 5767 12668 7380 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 9677 12699 9735 12705
rect 9677 12665 9689 12699
rect 9723 12696 9735 12699
rect 10778 12696 10784 12708
rect 9723 12668 10784 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 10778 12656 10784 12668
rect 10836 12656 10842 12708
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10134 12628 10140 12640
rect 10091 12600 10140 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 10505 12631 10563 12637
rect 10505 12597 10517 12631
rect 10551 12628 10563 12631
rect 11146 12628 11152 12640
rect 10551 12600 11152 12628
rect 10551 12597 10563 12600
rect 10505 12591 10563 12597
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 11330 12588 11336 12640
rect 11388 12588 11394 12640
rect 11793 12631 11851 12637
rect 11793 12597 11805 12631
rect 11839 12628 11851 12631
rect 11974 12628 11980 12640
rect 11839 12600 11980 12628
rect 11839 12597 11851 12600
rect 11793 12591 11851 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 1104 12538 12236 12560
rect 1104 12486 1550 12538
rect 1602 12486 1614 12538
rect 1666 12486 1678 12538
rect 1730 12486 1742 12538
rect 1794 12486 1806 12538
rect 1858 12486 3550 12538
rect 3602 12486 3614 12538
rect 3666 12486 3678 12538
rect 3730 12486 3742 12538
rect 3794 12486 3806 12538
rect 3858 12486 5550 12538
rect 5602 12486 5614 12538
rect 5666 12486 5678 12538
rect 5730 12486 5742 12538
rect 5794 12486 5806 12538
rect 5858 12486 7550 12538
rect 7602 12486 7614 12538
rect 7666 12486 7678 12538
rect 7730 12486 7742 12538
rect 7794 12486 7806 12538
rect 7858 12486 9550 12538
rect 9602 12486 9614 12538
rect 9666 12486 9678 12538
rect 9730 12486 9742 12538
rect 9794 12486 9806 12538
rect 9858 12486 11550 12538
rect 11602 12486 11614 12538
rect 11666 12486 11678 12538
rect 11730 12486 11742 12538
rect 11794 12486 11806 12538
rect 11858 12486 12236 12538
rect 1104 12464 12236 12486
rect 5442 12384 5448 12436
rect 5500 12384 5506 12436
rect 5902 12384 5908 12436
rect 5960 12384 5966 12436
rect 10045 12427 10103 12433
rect 10045 12393 10057 12427
rect 10091 12424 10103 12427
rect 12066 12424 12072 12436
rect 10091 12396 12072 12424
rect 10091 12393 10103 12396
rect 10045 12387 10103 12393
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 9861 12359 9919 12365
rect 9861 12325 9873 12359
rect 9907 12325 9919 12359
rect 9861 12319 9919 12325
rect 10321 12359 10379 12365
rect 10321 12325 10333 12359
rect 10367 12356 10379 12359
rect 10594 12356 10600 12368
rect 10367 12328 10600 12356
rect 10367 12325 10379 12328
rect 10321 12319 10379 12325
rect 5166 12248 5172 12300
rect 5224 12288 5230 12300
rect 6549 12291 6607 12297
rect 5224 12260 5580 12288
rect 5224 12248 5230 12260
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3936 12192 3985 12220
rect 3936 12180 3942 12192
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 4479 12192 4629 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 5552 12229 5580 12260
rect 6549 12257 6561 12291
rect 6595 12288 6607 12291
rect 6638 12288 6644 12300
rect 6595 12260 6644 12288
rect 6595 12257 6607 12260
rect 6549 12251 6607 12257
rect 6638 12248 6644 12260
rect 6696 12248 6702 12300
rect 9876 12288 9904 12319
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 10042 12288 10048 12300
rect 9876 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12288 10106 12300
rect 10873 12291 10931 12297
rect 10100 12260 10640 12288
rect 10100 12248 10106 12260
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 5316 12192 5365 12220
rect 5316 12180 5322 12192
rect 5353 12189 5365 12192
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12220 5595 12223
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 5583 12192 6837 12220
rect 5583 12189 5595 12192
rect 5537 12183 5595 12189
rect 6825 12189 6837 12192
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 5368 12152 5396 12183
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7101 12223 7159 12229
rect 7101 12220 7113 12223
rect 6972 12192 7113 12220
rect 6972 12180 6978 12192
rect 7101 12189 7113 12192
rect 7147 12189 7159 12223
rect 7101 12183 7159 12189
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 9364 12192 9413 12220
rect 9364 12180 9370 12192
rect 9401 12189 9413 12192
rect 9447 12220 9459 12223
rect 9950 12220 9956 12232
rect 9447 12192 9956 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10446 12223 10504 12229
rect 10446 12220 10458 12223
rect 10060 12192 10458 12220
rect 6641 12155 6699 12161
rect 6641 12152 6653 12155
rect 5368 12124 6653 12152
rect 6641 12121 6653 12124
rect 6687 12121 6699 12155
rect 6641 12115 6699 12121
rect 10060 12096 10088 12192
rect 10446 12189 10458 12192
rect 10492 12189 10504 12223
rect 10612 12220 10640 12260
rect 10873 12257 10885 12291
rect 10919 12288 10931 12291
rect 11149 12291 11207 12297
rect 11149 12288 11161 12291
rect 10919 12260 11161 12288
rect 10919 12257 10931 12260
rect 10873 12251 10931 12257
rect 11149 12257 11161 12260
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 10965 12223 11023 12229
rect 10965 12220 10977 12223
rect 10612 12192 10977 12220
rect 10446 12183 10504 12189
rect 10965 12189 10977 12192
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 11701 12223 11759 12229
rect 11701 12220 11713 12223
rect 11480 12192 11713 12220
rect 11480 12180 11486 12192
rect 11701 12189 11713 12192
rect 11747 12189 11759 12223
rect 11701 12183 11759 12189
rect 10229 12155 10287 12161
rect 10229 12121 10241 12155
rect 10275 12152 10287 12155
rect 10318 12152 10324 12164
rect 10275 12124 10324 12152
rect 10275 12121 10287 12124
rect 10229 12115 10287 12121
rect 10318 12112 10324 12124
rect 10376 12152 10382 12164
rect 10686 12152 10692 12164
rect 10376 12124 10692 12152
rect 10376 12112 10382 12124
rect 10686 12112 10692 12124
rect 10744 12112 10750 12164
rect 4062 12044 4068 12096
rect 4120 12044 4126 12096
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4341 12087 4399 12093
rect 4341 12084 4353 12087
rect 4212 12056 4353 12084
rect 4212 12044 4218 12056
rect 4341 12053 4353 12056
rect 4387 12053 4399 12087
rect 4341 12047 4399 12053
rect 5902 12044 5908 12096
rect 5960 12084 5966 12096
rect 7009 12087 7067 12093
rect 7009 12084 7021 12087
rect 5960 12056 7021 12084
rect 5960 12044 5966 12056
rect 7009 12053 7021 12056
rect 7055 12053 7067 12087
rect 7009 12047 7067 12053
rect 7190 12044 7196 12096
rect 7248 12044 7254 12096
rect 9490 12044 9496 12096
rect 9548 12044 9554 12096
rect 10042 12093 10048 12096
rect 10029 12087 10048 12093
rect 10029 12053 10041 12087
rect 10029 12047 10048 12053
rect 10042 12044 10048 12047
rect 10100 12044 10106 12096
rect 10505 12087 10563 12093
rect 10505 12053 10517 12087
rect 10551 12084 10563 12087
rect 12158 12084 12164 12096
rect 10551 12056 12164 12084
rect 10551 12053 10563 12056
rect 10505 12047 10563 12053
rect 12158 12044 12164 12056
rect 12216 12044 12222 12096
rect 1104 11994 12236 12016
rect 1104 11942 2250 11994
rect 2302 11942 2314 11994
rect 2366 11942 2378 11994
rect 2430 11942 2442 11994
rect 2494 11942 2506 11994
rect 2558 11942 4250 11994
rect 4302 11942 4314 11994
rect 4366 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 6250 11994
rect 6302 11942 6314 11994
rect 6366 11942 6378 11994
rect 6430 11942 6442 11994
rect 6494 11942 6506 11994
rect 6558 11942 8250 11994
rect 8302 11942 8314 11994
rect 8366 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 10250 11994
rect 10302 11942 10314 11994
rect 10366 11942 10378 11994
rect 10430 11942 10442 11994
rect 10494 11942 10506 11994
rect 10558 11942 12236 11994
rect 1104 11920 12236 11942
rect 4154 11880 4160 11892
rect 3344 11852 4160 11880
rect 3344 11821 3372 11852
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5442 11840 5448 11892
rect 5500 11840 5506 11892
rect 3329 11815 3387 11821
rect 3329 11781 3341 11815
rect 3375 11781 3387 11815
rect 3329 11775 3387 11781
rect 4062 11772 4068 11824
rect 4120 11772 4126 11824
rect 5460 11812 5488 11840
rect 5460 11784 5764 11812
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 3050 11636 3056 11688
rect 3108 11636 3114 11688
rect 5276 11676 5304 11707
rect 5350 11704 5356 11756
rect 5408 11704 5414 11756
rect 5442 11704 5448 11756
rect 5500 11704 5506 11756
rect 5736 11753 5764 11784
rect 7190 11772 7196 11824
rect 7248 11772 7254 11824
rect 9490 11772 9496 11824
rect 9548 11772 9554 11824
rect 10962 11772 10968 11824
rect 11020 11812 11026 11824
rect 11020 11784 11284 11812
rect 11020 11772 11026 11784
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10870 11744 10876 11756
rect 10100 11716 10876 11744
rect 10100 11704 10106 11716
rect 10870 11704 10876 11716
rect 10928 11744 10934 11756
rect 11057 11747 11115 11753
rect 11057 11744 11069 11747
rect 10928 11716 11069 11744
rect 10928 11704 10934 11716
rect 11057 11713 11069 11716
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11256 11744 11284 11784
rect 11330 11772 11336 11824
rect 11388 11772 11394 11824
rect 11609 11747 11667 11753
rect 11609 11744 11621 11747
rect 11256 11716 11621 11744
rect 11609 11713 11621 11716
rect 11655 11713 11667 11747
rect 11609 11707 11667 11713
rect 5994 11676 6000 11688
rect 5276 11648 6000 11676
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 7837 11679 7895 11685
rect 7837 11676 7849 11679
rect 7432 11648 7849 11676
rect 7432 11636 7438 11648
rect 7837 11645 7849 11648
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8481 11679 8539 11685
rect 8481 11676 8493 11679
rect 8159 11648 8493 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 8481 11645 8493 11648
rect 8527 11645 8539 11679
rect 8481 11639 8539 11645
rect 4801 11611 4859 11617
rect 4801 11577 4813 11611
rect 4847 11608 4859 11611
rect 5166 11608 5172 11620
rect 4847 11580 5172 11608
rect 4847 11577 4859 11580
rect 4801 11571 4859 11577
rect 5166 11568 5172 11580
rect 5224 11608 5230 11620
rect 5629 11611 5687 11617
rect 5629 11608 5641 11611
rect 5224 11580 5641 11608
rect 5224 11568 5230 11580
rect 5629 11577 5641 11580
rect 5675 11577 5687 11611
rect 6365 11611 6423 11617
rect 6365 11608 6377 11611
rect 5629 11571 5687 11577
rect 5920 11580 6377 11608
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 5077 11543 5135 11549
rect 5077 11540 5089 11543
rect 4028 11512 5089 11540
rect 4028 11500 4034 11512
rect 5077 11509 5089 11512
rect 5123 11509 5135 11543
rect 5077 11503 5135 11509
rect 5350 11500 5356 11552
rect 5408 11540 5414 11552
rect 5920 11540 5948 11580
rect 6365 11577 6377 11580
rect 6411 11608 6423 11611
rect 6638 11608 6644 11620
rect 6411 11580 6644 11608
rect 6411 11577 6423 11580
rect 6365 11571 6423 11577
rect 6638 11568 6644 11580
rect 6696 11568 6702 11620
rect 5408 11512 5948 11540
rect 5408 11500 5414 11512
rect 6086 11500 6092 11552
rect 6144 11500 6150 11552
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 8128 11540 8156 11639
rect 8754 11636 8760 11688
rect 8812 11636 8818 11688
rect 9214 11636 9220 11688
rect 9272 11676 9278 11688
rect 10060 11676 10088 11704
rect 9272 11648 10088 11676
rect 10229 11679 10287 11685
rect 9272 11636 9278 11648
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 10686 11676 10692 11688
rect 10275 11648 10692 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 10686 11636 10692 11648
rect 10744 11676 10750 11688
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 10744 11648 10977 11676
rect 10744 11636 10750 11648
rect 10965 11645 10977 11648
rect 11011 11676 11023 11679
rect 11164 11676 11192 11704
rect 11011 11648 11192 11676
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 10042 11568 10048 11620
rect 10100 11608 10106 11620
rect 10321 11611 10379 11617
rect 10321 11608 10333 11611
rect 10100 11580 10333 11608
rect 10100 11568 10106 11580
rect 10321 11577 10333 11580
rect 10367 11577 10379 11611
rect 10321 11571 10379 11577
rect 11238 11568 11244 11620
rect 11296 11608 11302 11620
rect 11333 11611 11391 11617
rect 11333 11608 11345 11611
rect 11296 11580 11345 11608
rect 11296 11568 11302 11580
rect 11333 11577 11345 11580
rect 11379 11577 11391 11611
rect 11333 11571 11391 11577
rect 9950 11540 9956 11552
rect 7156 11512 9956 11540
rect 7156 11500 7162 11512
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 11793 11543 11851 11549
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 11882 11540 11888 11552
rect 11839 11512 11888 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 1104 11450 12236 11472
rect 1104 11398 1550 11450
rect 1602 11398 1614 11450
rect 1666 11398 1678 11450
rect 1730 11398 1742 11450
rect 1794 11398 1806 11450
rect 1858 11398 3550 11450
rect 3602 11398 3614 11450
rect 3666 11398 3678 11450
rect 3730 11398 3742 11450
rect 3794 11398 3806 11450
rect 3858 11398 5550 11450
rect 5602 11398 5614 11450
rect 5666 11398 5678 11450
rect 5730 11398 5742 11450
rect 5794 11398 5806 11450
rect 5858 11398 7550 11450
rect 7602 11398 7614 11450
rect 7666 11398 7678 11450
rect 7730 11398 7742 11450
rect 7794 11398 7806 11450
rect 7858 11398 9550 11450
rect 9602 11398 9614 11450
rect 9666 11398 9678 11450
rect 9730 11398 9742 11450
rect 9794 11398 9806 11450
rect 9858 11398 11550 11450
rect 11602 11398 11614 11450
rect 11666 11398 11678 11450
rect 11730 11398 11742 11450
rect 11794 11398 11806 11450
rect 11858 11398 12236 11450
rect 1104 11376 12236 11398
rect 4617 11339 4675 11345
rect 4617 11336 4629 11339
rect 4356 11308 4629 11336
rect 4356 11277 4384 11308
rect 4617 11305 4629 11308
rect 4663 11305 4675 11339
rect 4617 11299 4675 11305
rect 5258 11296 5264 11348
rect 5316 11336 5322 11348
rect 5442 11336 5448 11348
rect 5316 11308 5448 11336
rect 5316 11296 5322 11308
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6914 11296 6920 11348
rect 6972 11296 6978 11348
rect 8754 11296 8760 11348
rect 8812 11336 8818 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8812 11308 8953 11336
rect 8812 11296 8818 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 11885 11339 11943 11345
rect 11885 11305 11897 11339
rect 11931 11336 11943 11339
rect 12066 11336 12072 11348
rect 11931 11308 12072 11336
rect 11931 11305 11943 11308
rect 11885 11299 11943 11305
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 4341 11271 4399 11277
rect 4341 11237 4353 11271
rect 4387 11237 4399 11271
rect 5350 11268 5356 11280
rect 4341 11231 4399 11237
rect 4816 11240 5356 11268
rect 3970 11160 3976 11212
rect 4028 11160 4034 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4614 11200 4620 11212
rect 4479 11172 4620 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 4816 11209 4844 11240
rect 5350 11228 5356 11240
rect 5408 11228 5414 11280
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11169 4859 11203
rect 4801 11163 4859 11169
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5994 11200 6000 11212
rect 5123 11172 6000 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6086 11160 6092 11212
rect 6144 11200 6150 11212
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 6144 11172 6745 11200
rect 6144 11160 6150 11172
rect 6733 11169 6745 11172
rect 6779 11169 6791 11203
rect 6932 11200 6960 11296
rect 10134 11228 10140 11280
rect 10192 11228 10198 11280
rect 6932 11172 7328 11200
rect 6733 11163 6791 11169
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11132 5043 11135
rect 5166 11132 5172 11144
rect 5031 11104 5172 11132
rect 5031 11101 5043 11104
rect 4985 11095 5043 11101
rect 4908 11064 4936 11095
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 7006 11092 7012 11144
rect 7064 11092 7070 11144
rect 7300 11141 7328 11172
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 9214 11200 9220 11212
rect 8628 11172 9220 11200
rect 8628 11160 8634 11172
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 10042 11200 10048 11212
rect 9324 11172 10048 11200
rect 9324 11141 9352 11172
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10152 11200 10180 11228
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 10152 11172 10425 11200
rect 10413 11169 10425 11172
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 10008 11104 10149 11132
rect 10008 11092 10014 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 5258 11064 5264 11076
rect 4908 11036 5264 11064
rect 5258 11024 5264 11036
rect 5316 11024 5322 11076
rect 7193 11067 7251 11073
rect 7193 11064 7205 11067
rect 6302 11036 6684 11064
rect 1946 10956 1952 11008
rect 2004 10996 2010 11008
rect 3970 10996 3976 11008
rect 2004 10968 3976 10996
rect 2004 10956 2010 10968
rect 3970 10956 3976 10968
rect 4028 10956 4034 11008
rect 6656 10996 6684 11036
rect 6840 11036 7205 11064
rect 6840 10996 6868 11036
rect 7193 11033 7205 11036
rect 7239 11033 7251 11067
rect 7193 11027 7251 11033
rect 11054 11024 11060 11076
rect 11112 11024 11118 11076
rect 6656 10968 6868 10996
rect 1104 10906 12236 10928
rect 1104 10854 2250 10906
rect 2302 10854 2314 10906
rect 2366 10854 2378 10906
rect 2430 10854 2442 10906
rect 2494 10854 2506 10906
rect 2558 10854 4250 10906
rect 4302 10854 4314 10906
rect 4366 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 6250 10906
rect 6302 10854 6314 10906
rect 6366 10854 6378 10906
rect 6430 10854 6442 10906
rect 6494 10854 6506 10906
rect 6558 10854 8250 10906
rect 8302 10854 8314 10906
rect 8366 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 10250 10906
rect 10302 10854 10314 10906
rect 10366 10854 10378 10906
rect 10430 10854 10442 10906
rect 10494 10854 10506 10906
rect 10558 10854 12236 10906
rect 1104 10832 12236 10854
rect 5629 10795 5687 10801
rect 5629 10761 5641 10795
rect 5675 10792 5687 10795
rect 5994 10792 6000 10804
rect 5675 10764 6000 10792
rect 5675 10761 5687 10764
rect 5629 10755 5687 10761
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 11333 10795 11391 10801
rect 11333 10761 11345 10795
rect 11379 10792 11391 10795
rect 11422 10792 11428 10804
rect 11379 10764 11428 10792
rect 11379 10761 11391 10764
rect 11333 10755 11391 10761
rect 11422 10752 11428 10764
rect 11480 10792 11486 10804
rect 11717 10795 11775 10801
rect 11717 10792 11729 10795
rect 11480 10764 11729 10792
rect 11480 10752 11486 10764
rect 11717 10761 11729 10764
rect 11763 10761 11775 10795
rect 11717 10755 11775 10761
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 12158 10792 12164 10804
rect 11931 10764 12164 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 3050 10684 3056 10736
rect 3108 10724 3114 10736
rect 4062 10724 4068 10736
rect 3108 10696 4068 10724
rect 3108 10684 3114 10696
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2682 10656 2688 10668
rect 1719 10628 2688 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3896 10665 3924 10696
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 4890 10684 4896 10736
rect 4948 10684 4954 10736
rect 9950 10724 9956 10736
rect 9600 10696 9956 10724
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 8754 10656 8760 10668
rect 8527 10628 8760 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9600 10665 9628 10696
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 11146 10684 11152 10736
rect 11204 10724 11210 10736
rect 11517 10727 11575 10733
rect 11517 10724 11529 10727
rect 11204 10696 11529 10724
rect 11204 10684 11210 10696
rect 11517 10693 11529 10696
rect 11563 10693 11575 10727
rect 11517 10687 11575 10693
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 9088 10628 9505 10656
rect 9088 10616 9094 10628
rect 9493 10625 9505 10628
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 4157 10591 4215 10597
rect 4157 10557 4169 10591
rect 4203 10588 4215 10591
rect 4614 10588 4620 10600
rect 4203 10560 4620 10588
rect 4203 10557 4215 10560
rect 4157 10551 4215 10557
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 8662 10548 8668 10600
rect 8720 10548 8726 10600
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10588 9919 10591
rect 10594 10588 10600 10600
rect 9907 10560 10600 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 10980 10588 11008 10642
rect 11054 10588 11060 10600
rect 10980 10560 11060 10588
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 12066 10520 12072 10532
rect 11716 10492 12072 10520
rect 842 10412 848 10464
rect 900 10452 906 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 900 10424 1501 10452
rect 900 10412 906 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 1489 10415 1547 10421
rect 8297 10455 8355 10461
rect 8297 10421 8309 10455
rect 8343 10452 8355 10455
rect 8570 10452 8576 10464
rect 8343 10424 8576 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 11716 10461 11744 10492
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9364 10424 9413 10452
rect 9364 10412 9370 10424
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 11701 10455 11759 10461
rect 11701 10421 11713 10455
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 1104 10362 12236 10384
rect 1104 10310 1550 10362
rect 1602 10310 1614 10362
rect 1666 10310 1678 10362
rect 1730 10310 1742 10362
rect 1794 10310 1806 10362
rect 1858 10310 3550 10362
rect 3602 10310 3614 10362
rect 3666 10310 3678 10362
rect 3730 10310 3742 10362
rect 3794 10310 3806 10362
rect 3858 10310 5550 10362
rect 5602 10310 5614 10362
rect 5666 10310 5678 10362
rect 5730 10310 5742 10362
rect 5794 10310 5806 10362
rect 5858 10310 7550 10362
rect 7602 10310 7614 10362
rect 7666 10310 7678 10362
rect 7730 10310 7742 10362
rect 7794 10310 7806 10362
rect 7858 10310 9550 10362
rect 9602 10310 9614 10362
rect 9666 10310 9678 10362
rect 9730 10310 9742 10362
rect 9794 10310 9806 10362
rect 9858 10310 11550 10362
rect 11602 10310 11614 10362
rect 11666 10310 11678 10362
rect 11730 10310 11742 10362
rect 11794 10310 11806 10362
rect 11858 10310 12236 10362
rect 1104 10288 12236 10310
rect 4890 10208 4896 10260
rect 4948 10208 4954 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11974 10248 11980 10260
rect 11655 10220 11980 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 1486 10072 1492 10124
rect 1544 10072 1550 10124
rect 1946 10072 1952 10124
rect 2004 10072 2010 10124
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 3145 10115 3203 10121
rect 3145 10112 3157 10115
rect 2740 10084 3157 10112
rect 2740 10072 2746 10084
rect 3145 10081 3157 10084
rect 3191 10081 3203 10115
rect 6914 10112 6920 10124
rect 3145 10075 3203 10081
rect 3896 10084 6920 10112
rect 3896 10056 3924 10084
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 2593 10047 2651 10053
rect 2593 10044 2605 10047
rect 1903 10016 2605 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 2593 10013 2605 10016
rect 2639 10013 2651 10047
rect 2593 10007 2651 10013
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10044 3571 10047
rect 3878 10044 3884 10056
rect 3559 10016 3884 10044
rect 3559 10013 3571 10016
rect 3513 10007 3571 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4614 10044 4620 10056
rect 4203 10016 4620 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 3326 9936 3332 9988
rect 3384 9976 3390 9988
rect 3789 9979 3847 9985
rect 3789 9976 3801 9979
rect 3384 9948 3801 9976
rect 3384 9936 3390 9948
rect 3789 9945 3801 9948
rect 3835 9945 3847 9979
rect 3988 9976 4016 10007
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 4816 10053 4844 10084
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 8846 10112 8852 10124
rect 8036 10084 8852 10112
rect 8036 10053 8064 10084
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 8297 10047 8355 10053
rect 8297 10013 8309 10047
rect 8343 10044 8355 10047
rect 8478 10044 8484 10056
rect 8343 10016 8484 10044
rect 8343 10013 8355 10016
rect 8297 10007 8355 10013
rect 5902 9976 5908 9988
rect 3988 9948 5908 9976
rect 3789 9939 3847 9945
rect 5902 9936 5908 9948
rect 5960 9936 5966 9988
rect 7852 9976 7880 10007
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 9766 10044 9772 10056
rect 8803 10016 9772 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 10962 10004 10968 10056
rect 11020 10004 11026 10056
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 8588 9976 8616 10004
rect 7852 9948 8616 9976
rect 8938 9936 8944 9988
rect 8996 9936 9002 9988
rect 11057 9979 11115 9985
rect 11057 9976 11069 9979
rect 9600 9948 11069 9976
rect 3418 9868 3424 9920
rect 3476 9868 3482 9920
rect 7282 9868 7288 9920
rect 7340 9908 7346 9920
rect 7929 9911 7987 9917
rect 7929 9908 7941 9911
rect 7340 9880 7941 9908
rect 7340 9868 7346 9880
rect 7929 9877 7941 9880
rect 7975 9877 7987 9911
rect 7929 9871 7987 9877
rect 8110 9868 8116 9920
rect 8168 9868 8174 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 9600 9908 9628 9948
rect 11057 9945 11069 9948
rect 11103 9976 11115 9979
rect 11238 9976 11244 9988
rect 11103 9948 11244 9976
rect 11103 9945 11115 9948
rect 11057 9939 11115 9945
rect 11238 9936 11244 9948
rect 11296 9936 11302 9988
rect 11330 9936 11336 9988
rect 11388 9936 11394 9988
rect 8720 9880 9628 9908
rect 8720 9868 8726 9880
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 10229 9911 10287 9917
rect 10229 9908 10241 9911
rect 10008 9880 10241 9908
rect 10008 9868 10014 9880
rect 10229 9877 10241 9880
rect 10275 9877 10287 9911
rect 10229 9871 10287 9877
rect 10778 9868 10784 9920
rect 10836 9868 10842 9920
rect 11149 9911 11207 9917
rect 11149 9877 11161 9911
rect 11195 9908 11207 9911
rect 11422 9908 11428 9920
rect 11195 9880 11428 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 1104 9818 12236 9840
rect 1104 9766 2250 9818
rect 2302 9766 2314 9818
rect 2366 9766 2378 9818
rect 2430 9766 2442 9818
rect 2494 9766 2506 9818
rect 2558 9766 4250 9818
rect 4302 9766 4314 9818
rect 4366 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 6250 9818
rect 6302 9766 6314 9818
rect 6366 9766 6378 9818
rect 6430 9766 6442 9818
rect 6494 9766 6506 9818
rect 6558 9766 8250 9818
rect 8302 9766 8314 9818
rect 8366 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 10250 9818
rect 10302 9766 10314 9818
rect 10366 9766 10378 9818
rect 10430 9766 10442 9818
rect 10494 9766 10506 9818
rect 10558 9766 12236 9818
rect 1104 9744 12236 9766
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 3237 9707 3295 9713
rect 3237 9704 3249 9707
rect 2740 9676 3249 9704
rect 2740 9664 2746 9676
rect 3237 9673 3249 9676
rect 3283 9704 3295 9707
rect 8938 9704 8944 9716
rect 3283 9676 4108 9704
rect 3283 9673 3295 9676
rect 3237 9667 3295 9673
rect 1486 9596 1492 9648
rect 1544 9636 1550 9648
rect 1765 9639 1823 9645
rect 1765 9636 1777 9639
rect 1544 9608 1777 9636
rect 1544 9596 1550 9608
rect 1765 9605 1777 9608
rect 1811 9605 1823 9639
rect 3418 9636 3424 9648
rect 2990 9608 3424 9636
rect 1765 9599 1823 9605
rect 3418 9596 3424 9608
rect 3476 9596 3482 9648
rect 4080 9636 4108 9676
rect 8312 9676 8944 9704
rect 5442 9636 5448 9648
rect 4080 9608 5448 9636
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 5537 9639 5595 9645
rect 5537 9605 5549 9639
rect 5583 9636 5595 9639
rect 6638 9636 6644 9648
rect 5583 9608 6644 9636
rect 5583 9605 5595 9608
rect 5537 9599 5595 9605
rect 6638 9596 6644 9608
rect 6696 9636 6702 9648
rect 8312 9636 8340 9676
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 6696 9608 8340 9636
rect 6696 9596 6702 9608
rect 9766 9596 9772 9648
rect 9824 9596 9830 9648
rect 10042 9596 10048 9648
rect 10100 9636 10106 9648
rect 10870 9636 10876 9648
rect 10100 9608 10876 9636
rect 10100 9596 10106 9608
rect 10870 9596 10876 9608
rect 10928 9636 10934 9648
rect 11701 9639 11759 9645
rect 11701 9636 11713 9639
rect 10928 9608 11713 9636
rect 10928 9596 10934 9608
rect 11701 9605 11713 9608
rect 11747 9605 11759 9639
rect 11701 9599 11759 9605
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 7650 9568 7656 9580
rect 6972 9540 7656 9568
rect 6972 9528 6978 9540
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 9692 9540 10425 9568
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 1489 9503 1547 9509
rect 1489 9500 1501 9503
rect 1452 9472 1501 9500
rect 1452 9460 1458 9472
rect 1489 9469 1501 9472
rect 1535 9469 1547 9503
rect 1489 9463 1547 9469
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 7929 9503 7987 9509
rect 7929 9500 7941 9503
rect 7064 9472 7941 9500
rect 7064 9460 7070 9472
rect 7929 9469 7941 9472
rect 7975 9469 7987 9503
rect 7929 9463 7987 9469
rect 8202 9460 8208 9512
rect 8260 9460 8266 9512
rect 9692 9509 9720 9540
rect 10413 9537 10425 9540
rect 10459 9568 10471 9571
rect 10962 9568 10968 9580
rect 10459 9540 10968 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11379 9540 11529 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9568 11851 9571
rect 12158 9568 12164 9580
rect 11839 9540 12164 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9469 9735 9503
rect 9677 9463 9735 9469
rect 10781 9503 10839 9509
rect 10781 9469 10793 9503
rect 10827 9500 10839 9503
rect 11146 9500 11152 9512
rect 10827 9472 11152 9500
rect 10827 9469 10839 9472
rect 10781 9463 10839 9469
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 9398 9392 9404 9444
rect 9456 9432 9462 9444
rect 11517 9435 11575 9441
rect 11517 9432 11529 9435
rect 9456 9404 11529 9432
rect 9456 9392 9462 9404
rect 11517 9401 11529 9404
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 3970 9364 3976 9376
rect 2188 9336 3976 9364
rect 2188 9324 2194 9336
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4062 9324 4068 9376
rect 4120 9324 4126 9376
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 6086 9364 6092 9376
rect 4672 9336 6092 9364
rect 4672 9324 4678 9336
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 7745 9367 7803 9373
rect 7745 9333 7757 9367
rect 7791 9364 7803 9367
rect 7926 9364 7932 9376
rect 7791 9336 7932 9364
rect 7791 9333 7803 9336
rect 7745 9327 7803 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 1104 9274 12236 9296
rect 1104 9222 1550 9274
rect 1602 9222 1614 9274
rect 1666 9222 1678 9274
rect 1730 9222 1742 9274
rect 1794 9222 1806 9274
rect 1858 9222 3550 9274
rect 3602 9222 3614 9274
rect 3666 9222 3678 9274
rect 3730 9222 3742 9274
rect 3794 9222 3806 9274
rect 3858 9222 5550 9274
rect 5602 9222 5614 9274
rect 5666 9222 5678 9274
rect 5730 9222 5742 9274
rect 5794 9222 5806 9274
rect 5858 9222 7550 9274
rect 7602 9222 7614 9274
rect 7666 9222 7678 9274
rect 7730 9222 7742 9274
rect 7794 9222 7806 9274
rect 7858 9222 9550 9274
rect 9602 9222 9614 9274
rect 9666 9222 9678 9274
rect 9730 9222 9742 9274
rect 9794 9222 9806 9274
rect 9858 9222 11550 9274
rect 11602 9222 11614 9274
rect 11666 9222 11678 9274
rect 11730 9222 11742 9274
rect 11794 9222 11806 9274
rect 11858 9222 12236 9274
rect 1104 9200 12236 9222
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 5537 9163 5595 9169
rect 2924 9132 3556 9160
rect 2924 9120 2930 9132
rect 842 9052 848 9104
rect 900 9092 906 9104
rect 1489 9095 1547 9101
rect 1489 9092 1501 9095
rect 900 9064 1501 9092
rect 900 9052 906 9064
rect 1489 9061 1501 9064
rect 1535 9061 1547 9095
rect 1489 9055 1547 9061
rect 1857 9095 1915 9101
rect 1857 9061 1869 9095
rect 1903 9092 1915 9095
rect 2130 9092 2136 9104
rect 1903 9064 2136 9092
rect 1903 9061 1915 9064
rect 1857 9055 1915 9061
rect 2130 9052 2136 9064
rect 2188 9052 2194 9104
rect 3528 9092 3556 9132
rect 5537 9129 5549 9163
rect 5583 9160 5595 9163
rect 5902 9160 5908 9172
rect 5583 9132 5908 9160
rect 5583 9129 5595 9132
rect 5537 9123 5595 9129
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 6086 9120 6092 9172
rect 6144 9120 6150 9172
rect 8662 9120 8668 9172
rect 8720 9160 8726 9172
rect 8757 9163 8815 9169
rect 8757 9160 8769 9163
rect 8720 9132 8769 9160
rect 8720 9120 8726 9132
rect 8757 9129 8769 9132
rect 8803 9129 8815 9163
rect 8757 9123 8815 9129
rect 6549 9095 6607 9101
rect 6549 9092 6561 9095
rect 3528 9064 6561 9092
rect 6549 9061 6561 9064
rect 6595 9061 6607 9095
rect 6549 9055 6607 9061
rect 1394 8984 1400 9036
rect 1452 9024 1458 9036
rect 3605 9027 3663 9033
rect 3605 9024 3617 9027
rect 1452 8996 3617 9024
rect 1452 8984 1458 8996
rect 3605 8993 3617 8996
rect 3651 9024 3663 9027
rect 4062 9024 4068 9036
rect 3651 8996 4068 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 3804 8968 3832 8996
rect 4062 8984 4068 8996
rect 4120 9024 4126 9036
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 4120 8996 7021 9024
rect 4120 8984 4126 8996
rect 7009 8993 7021 8996
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 7282 8984 7288 9036
rect 7340 8984 7346 9036
rect 8772 9024 8800 9123
rect 10042 9120 10048 9172
rect 10100 9120 10106 9172
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 8772 8996 9505 9024
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10137 9027 10195 9033
rect 10137 9024 10149 9027
rect 10008 8996 10149 9024
rect 10008 8984 10014 8996
rect 10137 8993 10149 8996
rect 10183 8993 10195 9027
rect 10137 8987 10195 8993
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 2038 8956 2044 8968
rect 1719 8928 2044 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 3786 8916 3792 8968
rect 3844 8916 3850 8968
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4028 8928 5304 8956
rect 4028 8916 4034 8928
rect 2866 8848 2872 8900
rect 2924 8848 2930 8900
rect 3326 8848 3332 8900
rect 3384 8848 3390 8900
rect 3418 8848 3424 8900
rect 3476 8888 3482 8900
rect 4614 8888 4620 8900
rect 3476 8860 4620 8888
rect 3476 8848 3482 8860
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 5276 8888 5304 8928
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 5721 8959 5779 8965
rect 5721 8958 5733 8959
rect 5644 8930 5733 8958
rect 5644 8888 5672 8930
rect 5721 8925 5733 8930
rect 5767 8958 5779 8959
rect 5767 8956 5856 8958
rect 5902 8956 5908 8968
rect 5767 8930 5908 8956
rect 5767 8925 5779 8930
rect 5828 8928 5908 8930
rect 5721 8919 5779 8925
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 5994 8916 6000 8968
rect 6052 8916 6058 8968
rect 6086 8916 6092 8968
rect 6144 8916 6150 8968
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 6730 8956 6736 8968
rect 6687 8928 6736 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 8864 8928 9781 8956
rect 5276 8860 5672 8888
rect 6178 8848 6184 8900
rect 6236 8848 6242 8900
rect 6365 8891 6423 8897
rect 6365 8857 6377 8891
rect 6411 8857 6423 8891
rect 6365 8851 6423 8857
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 3292 8792 4813 8820
rect 3292 8780 3298 8792
rect 4801 8789 4813 8792
rect 4847 8789 4859 8823
rect 4801 8783 4859 8789
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 5905 8823 5963 8829
rect 5905 8820 5917 8823
rect 5500 8792 5917 8820
rect 5500 8780 5506 8792
rect 5905 8789 5917 8792
rect 5951 8789 5963 8823
rect 5905 8783 5963 8789
rect 5994 8780 6000 8832
rect 6052 8820 6058 8832
rect 6380 8820 6408 8851
rect 7926 8848 7932 8900
rect 7984 8848 7990 8900
rect 6052 8792 6408 8820
rect 6052 8780 6058 8792
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 8864 8820 8892 8928
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 10042 8956 10048 8968
rect 9907 8928 10048 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9490 8888 9496 8900
rect 9088 8860 9496 8888
rect 9088 8848 9094 8860
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 8076 8792 8892 8820
rect 8941 8823 8999 8829
rect 8076 8780 8082 8792
rect 8941 8789 8953 8823
rect 8987 8820 8999 8823
rect 9122 8820 9128 8832
rect 8987 8792 9128 8820
rect 8987 8789 8999 8792
rect 8941 8783 8999 8789
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9784 8820 9812 8919
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10413 8891 10471 8897
rect 10413 8888 10425 8891
rect 10008 8860 10425 8888
rect 10008 8848 10014 8860
rect 10413 8857 10425 8860
rect 10459 8857 10471 8891
rect 10413 8851 10471 8857
rect 10870 8848 10876 8900
rect 10928 8848 10934 8900
rect 9858 8820 9864 8832
rect 9784 8792 9864 8820
rect 9858 8780 9864 8792
rect 9916 8820 9922 8832
rect 10686 8820 10692 8832
rect 9916 8792 10692 8820
rect 9916 8780 9922 8792
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11204 8792 11897 8820
rect 11204 8780 11210 8792
rect 11885 8789 11897 8792
rect 11931 8789 11943 8823
rect 11885 8783 11943 8789
rect 1104 8730 12236 8752
rect 1104 8678 2250 8730
rect 2302 8678 2314 8730
rect 2366 8678 2378 8730
rect 2430 8678 2442 8730
rect 2494 8678 2506 8730
rect 2558 8678 4250 8730
rect 4302 8678 4314 8730
rect 4366 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 6250 8730
rect 6302 8678 6314 8730
rect 6366 8678 6378 8730
rect 6430 8678 6442 8730
rect 6494 8678 6506 8730
rect 6558 8678 8250 8730
rect 8302 8678 8314 8730
rect 8366 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 10250 8730
rect 10302 8678 10314 8730
rect 10366 8678 10378 8730
rect 10430 8678 10442 8730
rect 10494 8678 10506 8730
rect 10558 8678 12236 8730
rect 1104 8656 12236 8678
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 2225 8619 2283 8625
rect 2225 8616 2237 8619
rect 2188 8588 2237 8616
rect 2188 8576 2194 8588
rect 2225 8585 2237 8588
rect 2271 8585 2283 8619
rect 2225 8579 2283 8585
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 2590 8616 2596 8628
rect 2464 8588 2596 8616
rect 2464 8576 2470 8588
rect 2590 8576 2596 8588
rect 2648 8616 2654 8628
rect 5350 8616 5356 8628
rect 2648 8588 5356 8616
rect 2648 8576 2654 8588
rect 5350 8576 5356 8588
rect 5408 8616 5414 8628
rect 5537 8619 5595 8625
rect 5537 8616 5549 8619
rect 5408 8588 5549 8616
rect 5408 8576 5414 8588
rect 5537 8585 5549 8588
rect 5583 8585 5595 8619
rect 5537 8579 5595 8585
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8662 8616 8668 8628
rect 7975 8588 8668 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 8662 8576 8668 8588
rect 8720 8616 8726 8628
rect 9582 8616 9588 8628
rect 8720 8588 9588 8616
rect 8720 8576 8726 8588
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9769 8619 9827 8625
rect 9769 8585 9781 8619
rect 9815 8585 9827 8619
rect 9769 8579 9827 8585
rect 1946 8508 1952 8560
rect 2004 8548 2010 8560
rect 3326 8548 3332 8560
rect 2004 8520 3332 8548
rect 2004 8508 2010 8520
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2406 8480 2412 8492
rect 1719 8452 2412 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 2516 8489 2544 8520
rect 3326 8508 3332 8520
rect 3384 8508 3390 8560
rect 5721 8551 5779 8557
rect 5721 8548 5733 8551
rect 5290 8520 5733 8548
rect 5721 8517 5733 8520
rect 5767 8517 5779 8551
rect 8754 8548 8760 8560
rect 5721 8511 5779 8517
rect 7576 8520 8760 8548
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3786 8440 3792 8492
rect 3844 8440 3850 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6730 8480 6736 8492
rect 5859 8452 6736 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7576 8489 7604 8520
rect 8754 8508 8760 8520
rect 8812 8548 8818 8560
rect 9784 8548 9812 8579
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10100 8588 10609 8616
rect 10100 8576 10106 8588
rect 10597 8585 10609 8588
rect 10643 8616 10655 8619
rect 10778 8616 10784 8628
rect 10643 8588 10784 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 11793 8619 11851 8625
rect 11296 8588 11652 8616
rect 11296 8576 11302 8588
rect 8812 8520 9812 8548
rect 8812 8508 8818 8520
rect 9858 8508 9864 8560
rect 9916 8557 9922 8560
rect 9916 8551 9979 8557
rect 9916 8517 9933 8551
rect 9967 8517 9979 8551
rect 9916 8511 9979 8517
rect 9916 8508 9922 8511
rect 10134 8508 10140 8560
rect 10192 8508 10198 8560
rect 10873 8551 10931 8557
rect 10244 8520 10808 8548
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8480 7895 8483
rect 7926 8480 7932 8492
rect 7883 8452 7932 8480
rect 7883 8449 7895 8452
rect 7837 8443 7895 8449
rect 2038 8372 2044 8424
rect 2096 8372 2102 8424
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8412 2191 8415
rect 2314 8412 2320 8424
rect 2179 8384 2320 8412
rect 2179 8381 2191 8384
rect 2133 8375 2191 8381
rect 2314 8372 2320 8384
rect 2372 8412 2378 8424
rect 2682 8412 2688 8424
rect 2372 8384 2688 8412
rect 2372 8372 2378 8384
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3418 8412 3424 8424
rect 3375 8384 3424 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 3620 8384 4077 8412
rect 842 8304 848 8356
rect 900 8344 906 8356
rect 1489 8347 1547 8353
rect 1489 8344 1501 8347
rect 900 8316 1501 8344
rect 900 8304 906 8316
rect 1489 8313 1501 8316
rect 1535 8313 1547 8347
rect 1489 8307 1547 8313
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 1946 8344 1952 8356
rect 1903 8316 1952 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 1946 8304 1952 8316
rect 2004 8304 2010 8356
rect 3620 8353 3648 8384
rect 4065 8381 4077 8384
rect 4111 8381 4123 8415
rect 7760 8412 7788 8443
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 8159 8452 8493 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 9214 8440 9220 8492
rect 9272 8440 9278 8492
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 10152 8480 10180 8508
rect 9640 8452 10180 8480
rect 9640 8440 9646 8452
rect 7760 8384 8156 8412
rect 4065 8375 4123 8381
rect 8128 8353 8156 8384
rect 9030 8372 9036 8424
rect 9088 8372 9094 8424
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 10042 8412 10048 8424
rect 9548 8384 10048 8412
rect 9548 8372 9554 8384
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10244 8412 10272 8520
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 10152 8384 10272 8412
rect 10520 8412 10548 8443
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 10780 8480 10808 8520
rect 10873 8517 10885 8551
rect 10919 8548 10931 8551
rect 11146 8548 11152 8560
rect 10919 8520 11152 8548
rect 10919 8517 10931 8520
rect 10873 8511 10931 8517
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10780 8452 11069 8480
rect 11057 8449 11069 8452
rect 11103 8480 11115 8483
rect 11422 8480 11428 8492
rect 11103 8452 11428 8480
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 11624 8489 11652 8588
rect 11793 8585 11805 8619
rect 11839 8616 11851 8619
rect 12066 8616 12072 8628
rect 11839 8588 12072 8616
rect 11839 8585 11851 8588
rect 11793 8579 11851 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8449 11667 8483
rect 11609 8443 11667 8449
rect 12158 8412 12164 8424
rect 10520 8384 12164 8412
rect 3605 8347 3663 8353
rect 3605 8313 3617 8347
rect 3651 8313 3663 8347
rect 3605 8307 3663 8313
rect 8113 8347 8171 8353
rect 8113 8313 8125 8347
rect 8159 8313 8171 8347
rect 8113 8307 8171 8313
rect 9582 8304 9588 8356
rect 9640 8344 9646 8356
rect 10152 8344 10180 8384
rect 12158 8372 12164 8384
rect 12216 8372 12222 8424
rect 9640 8316 10180 8344
rect 9640 8304 9646 8316
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 5994 8276 6000 8288
rect 3384 8248 6000 8276
rect 3384 8236 3390 8248
rect 5994 8236 6000 8248
rect 6052 8236 6058 8288
rect 7282 8236 7288 8288
rect 7340 8276 7346 8288
rect 7561 8279 7619 8285
rect 7561 8276 7573 8279
rect 7340 8248 7573 8276
rect 7340 8236 7346 8248
rect 7561 8245 7573 8248
rect 7607 8245 7619 8279
rect 7561 8239 7619 8245
rect 9953 8279 10011 8285
rect 9953 8245 9965 8279
rect 9999 8276 10011 8279
rect 10152 8276 10180 8316
rect 11241 8347 11299 8353
rect 11241 8313 11253 8347
rect 11287 8344 11299 8347
rect 12066 8344 12072 8356
rect 11287 8316 12072 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 9999 8248 10180 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10318 8236 10324 8288
rect 10376 8236 10382 8288
rect 1104 8186 12236 8208
rect 1104 8134 1550 8186
rect 1602 8134 1614 8186
rect 1666 8134 1678 8186
rect 1730 8134 1742 8186
rect 1794 8134 1806 8186
rect 1858 8134 3550 8186
rect 3602 8134 3614 8186
rect 3666 8134 3678 8186
rect 3730 8134 3742 8186
rect 3794 8134 3806 8186
rect 3858 8134 5550 8186
rect 5602 8134 5614 8186
rect 5666 8134 5678 8186
rect 5730 8134 5742 8186
rect 5794 8134 5806 8186
rect 5858 8134 7550 8186
rect 7602 8134 7614 8186
rect 7666 8134 7678 8186
rect 7730 8134 7742 8186
rect 7794 8134 7806 8186
rect 7858 8134 9550 8186
rect 9602 8134 9614 8186
rect 9666 8134 9678 8186
rect 9730 8134 9742 8186
rect 9794 8134 9806 8186
rect 9858 8134 11550 8186
rect 11602 8134 11614 8186
rect 11666 8134 11678 8186
rect 11730 8134 11742 8186
rect 11794 8134 11806 8186
rect 11858 8134 12236 8186
rect 1104 8112 12236 8134
rect 6638 8032 6644 8084
rect 6696 8032 6702 8084
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8904 8044 8953 8072
rect 8904 8032 8910 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 9401 8075 9459 8081
rect 9401 8041 9413 8075
rect 9447 8072 9459 8075
rect 9950 8072 9956 8084
rect 9447 8044 9956 8072
rect 9447 8041 9459 8044
rect 9401 8035 9459 8041
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10781 8075 10839 8081
rect 10781 8041 10793 8075
rect 10827 8072 10839 8075
rect 10870 8072 10876 8084
rect 10827 8044 10876 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11054 8032 11060 8084
rect 11112 8032 11118 8084
rect 11793 8075 11851 8081
rect 11793 8041 11805 8075
rect 11839 8072 11851 8075
rect 11882 8072 11888 8084
rect 11839 8044 11888 8072
rect 11839 8041 11851 8044
rect 11793 8035 11851 8041
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 2314 7964 2320 8016
rect 2372 7964 2378 8016
rect 8757 8007 8815 8013
rect 8757 7973 8769 8007
rect 8803 8004 8815 8007
rect 9030 8004 9036 8016
rect 8803 7976 9036 8004
rect 8803 7973 8815 7976
rect 8757 7967 8815 7973
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 9214 7964 9220 8016
rect 9272 8004 9278 8016
rect 9272 7976 10732 8004
rect 9272 7964 9278 7976
rect 7282 7896 7288 7948
rect 7340 7896 7346 7948
rect 9950 7936 9956 7948
rect 9416 7908 9956 7936
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2038 7868 2044 7880
rect 1719 7840 2044 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2038 7828 2044 7840
rect 2096 7868 2102 7880
rect 2096 7840 2728 7868
rect 2096 7828 2102 7840
rect 2130 7760 2136 7812
rect 2188 7800 2194 7812
rect 2501 7803 2559 7809
rect 2501 7800 2513 7803
rect 2188 7772 2513 7800
rect 2188 7760 2194 7772
rect 2501 7769 2513 7772
rect 2547 7769 2559 7803
rect 2501 7763 2559 7769
rect 2590 7760 2596 7812
rect 2648 7760 2654 7812
rect 2700 7744 2728 7840
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4212 7840 5181 7868
rect 4212 7828 4218 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 7006 7828 7012 7880
rect 7064 7828 7070 7880
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8812 7840 8953 7868
rect 8812 7828 8818 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9122 7828 9128 7880
rect 9180 7828 9186 7880
rect 9416 7877 9444 7908
rect 9950 7896 9956 7908
rect 10008 7936 10014 7948
rect 10318 7936 10324 7948
rect 10008 7908 10324 7936
rect 10008 7896 10014 7908
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9548 7840 9597 7868
rect 9548 7828 9554 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 10042 7868 10048 7880
rect 9723 7840 10048 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10704 7877 10732 7976
rect 11146 7964 11152 8016
rect 11204 7964 11210 8016
rect 11164 7936 11192 7964
rect 11164 7908 11652 7936
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 11146 7868 11152 7880
rect 10735 7840 11152 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7868 11299 7871
rect 11330 7868 11336 7880
rect 11287 7840 11336 7868
rect 11287 7837 11299 7840
rect 11241 7831 11299 7837
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 11624 7877 11652 7908
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 9769 7803 9827 7809
rect 9769 7800 9781 7803
rect 8510 7772 9781 7800
rect 9769 7769 9781 7772
rect 9815 7769 9827 7803
rect 9769 7763 9827 7769
rect 842 7692 848 7744
rect 900 7732 906 7744
rect 1489 7735 1547 7741
rect 1489 7732 1501 7735
rect 900 7704 1501 7732
rect 900 7692 906 7704
rect 1489 7701 1501 7704
rect 1535 7701 1547 7735
rect 1489 7695 1547 7701
rect 2682 7692 2688 7744
rect 2740 7692 2746 7744
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 3418 7732 3424 7744
rect 2915 7704 3424 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 11422 7692 11428 7744
rect 11480 7692 11486 7744
rect 1104 7642 12236 7664
rect 1104 7590 2250 7642
rect 2302 7590 2314 7642
rect 2366 7590 2378 7642
rect 2430 7590 2442 7642
rect 2494 7590 2506 7642
rect 2558 7590 4250 7642
rect 4302 7590 4314 7642
rect 4366 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 6250 7642
rect 6302 7590 6314 7642
rect 6366 7590 6378 7642
rect 6430 7590 6442 7642
rect 6494 7590 6506 7642
rect 6558 7590 8250 7642
rect 8302 7590 8314 7642
rect 8366 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 10250 7642
rect 10302 7590 10314 7642
rect 10366 7590 10378 7642
rect 10430 7590 10442 7642
rect 10494 7590 10506 7642
rect 10558 7590 12236 7642
rect 1104 7568 12236 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3237 7531 3295 7537
rect 3237 7528 3249 7531
rect 2740 7500 3249 7528
rect 2740 7488 2746 7500
rect 3237 7497 3249 7500
rect 3283 7497 3295 7531
rect 3237 7491 3295 7497
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 8720 7500 8769 7528
rect 8720 7488 8726 7500
rect 8757 7497 8769 7500
rect 8803 7497 8815 7531
rect 8757 7491 8815 7497
rect 3421 7463 3479 7469
rect 3421 7460 3433 7463
rect 2990 7432 3433 7460
rect 3421 7429 3433 7432
rect 3467 7429 3479 7463
rect 9677 7463 9735 7469
rect 9677 7460 9689 7463
rect 8510 7432 9689 7460
rect 3421 7423 3479 7429
rect 9677 7429 9689 7432
rect 9723 7429 9735 7463
rect 9677 7423 9735 7429
rect 1394 7352 1400 7404
rect 1452 7392 1458 7404
rect 1489 7395 1547 7401
rect 1489 7392 1501 7395
rect 1452 7364 1501 7392
rect 1452 7352 1458 7364
rect 1489 7361 1501 7364
rect 1535 7361 1547 7395
rect 1489 7355 1547 7361
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3970 7392 3976 7404
rect 3559 7364 3976 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 8662 7352 8668 7404
rect 8720 7392 8726 7404
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 8720 7364 9413 7392
rect 8720 7352 8726 7364
rect 9401 7361 9413 7364
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7392 10471 7395
rect 10962 7392 10968 7404
rect 10459 7364 10968 7392
rect 10459 7361 10471 7364
rect 10413 7355 10471 7361
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 1854 7324 1860 7336
rect 1811 7296 1860 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 7282 7284 7288 7336
rect 7340 7284 7346 7336
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 9600 7324 9628 7355
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7392 11575 7395
rect 11563 7364 11597 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 9088 7296 9628 7324
rect 10781 7327 10839 7333
rect 9088 7284 9094 7296
rect 10781 7293 10793 7327
rect 10827 7324 10839 7327
rect 11532 7324 11560 7355
rect 11974 7324 11980 7336
rect 10827 7296 11980 7324
rect 10827 7293 10839 7296
rect 10781 7287 10839 7293
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 8294 7216 8300 7268
rect 8352 7256 8358 7268
rect 8849 7259 8907 7265
rect 8849 7256 8861 7259
rect 8352 7228 8861 7256
rect 8352 7216 8358 7228
rect 8849 7225 8861 7228
rect 8895 7225 8907 7259
rect 8849 7219 8907 7225
rect 10505 7191 10563 7197
rect 10505 7157 10517 7191
rect 10551 7188 10563 7191
rect 11238 7188 11244 7200
rect 10551 7160 11244 7188
rect 10551 7157 10563 7160
rect 10505 7151 10563 7157
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 11330 7148 11336 7200
rect 11388 7148 11394 7200
rect 11701 7191 11759 7197
rect 11701 7157 11713 7191
rect 11747 7188 11759 7191
rect 11882 7188 11888 7200
rect 11747 7160 11888 7188
rect 11747 7157 11759 7160
rect 11701 7151 11759 7157
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 1104 7098 12236 7120
rect 1104 7046 1550 7098
rect 1602 7046 1614 7098
rect 1666 7046 1678 7098
rect 1730 7046 1742 7098
rect 1794 7046 1806 7098
rect 1858 7046 3550 7098
rect 3602 7046 3614 7098
rect 3666 7046 3678 7098
rect 3730 7046 3742 7098
rect 3794 7046 3806 7098
rect 3858 7046 5550 7098
rect 5602 7046 5614 7098
rect 5666 7046 5678 7098
rect 5730 7046 5742 7098
rect 5794 7046 5806 7098
rect 5858 7046 7550 7098
rect 7602 7046 7614 7098
rect 7666 7046 7678 7098
rect 7730 7046 7742 7098
rect 7794 7046 7806 7098
rect 7858 7046 9550 7098
rect 9602 7046 9614 7098
rect 9666 7046 9678 7098
rect 9730 7046 9742 7098
rect 9794 7046 9806 7098
rect 9858 7046 11550 7098
rect 11602 7046 11614 7098
rect 11666 7046 11678 7098
rect 11730 7046 11742 7098
rect 11794 7046 11806 7098
rect 11858 7046 12236 7098
rect 1104 7024 12236 7046
rect 1765 6987 1823 6993
rect 1765 6953 1777 6987
rect 1811 6984 1823 6987
rect 1946 6984 1952 6996
rect 1811 6956 1952 6984
rect 1811 6953 1823 6956
rect 1765 6947 1823 6953
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 7101 6987 7159 6993
rect 7101 6953 7113 6987
rect 7147 6984 7159 6987
rect 7282 6984 7288 6996
rect 7147 6956 7288 6984
rect 7147 6953 7159 6956
rect 7101 6947 7159 6953
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 1857 6919 1915 6925
rect 1857 6885 1869 6919
rect 1903 6914 1915 6919
rect 9950 6916 9956 6928
rect 1903 6886 1937 6914
rect 9416 6888 9956 6916
rect 1903 6885 1915 6886
rect 1857 6879 1915 6885
rect 1872 6848 1900 6879
rect 2038 6848 2044 6860
rect 1872 6820 2044 6848
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7377 6851 7435 6857
rect 7377 6848 7389 6851
rect 6972 6820 7389 6848
rect 6972 6808 6978 6820
rect 7377 6817 7389 6820
rect 7423 6848 7435 6851
rect 7926 6848 7932 6860
rect 7423 6820 7932 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 8938 6808 8944 6860
rect 8996 6808 9002 6860
rect 9416 6857 9444 6888
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 9401 6851 9459 6857
rect 9401 6817 9413 6851
rect 9447 6817 9459 6851
rect 9968 6848 9996 6876
rect 10778 6848 10784 6860
rect 9968 6820 10784 6848
rect 9401 6811 9459 6817
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 7469 6783 7527 6789
rect 7469 6749 7481 6783
rect 7515 6780 7527 6783
rect 8294 6780 8300 6792
rect 7515 6752 8300 6780
rect 7515 6749 7527 6752
rect 7469 6743 7527 6749
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 8904 6752 9321 6780
rect 8904 6740 8910 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 2038 6672 2044 6724
rect 2096 6712 2102 6724
rect 2225 6715 2283 6721
rect 2225 6712 2237 6715
rect 2096 6684 2237 6712
rect 2096 6672 2102 6684
rect 2225 6681 2237 6684
rect 2271 6681 2283 6715
rect 2225 6675 2283 6681
rect 10134 6672 10140 6724
rect 10192 6712 10198 6724
rect 10229 6715 10287 6721
rect 10229 6712 10241 6715
rect 10192 6684 10241 6712
rect 10192 6672 10198 6684
rect 10229 6681 10241 6684
rect 10275 6681 10287 6715
rect 10229 6675 10287 6681
rect 11238 6672 11244 6724
rect 11296 6672 11302 6724
rect 11701 6647 11759 6653
rect 11701 6613 11713 6647
rect 11747 6644 11759 6647
rect 11974 6644 11980 6656
rect 11747 6616 11980 6644
rect 11747 6613 11759 6616
rect 11701 6607 11759 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 1104 6554 12236 6576
rect 1104 6502 2250 6554
rect 2302 6502 2314 6554
rect 2366 6502 2378 6554
rect 2430 6502 2442 6554
rect 2494 6502 2506 6554
rect 2558 6502 4250 6554
rect 4302 6502 4314 6554
rect 4366 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 6250 6554
rect 6302 6502 6314 6554
rect 6366 6502 6378 6554
rect 6430 6502 6442 6554
rect 6494 6502 6506 6554
rect 6558 6502 8250 6554
rect 8302 6502 8314 6554
rect 8366 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 10250 6554
rect 10302 6502 10314 6554
rect 10366 6502 10378 6554
rect 10430 6502 10442 6554
rect 10494 6502 10506 6554
rect 10558 6502 12236 6554
rect 1104 6480 12236 6502
rect 8846 6400 8852 6452
rect 8904 6400 8910 6452
rect 1946 6332 1952 6384
rect 2004 6332 2010 6384
rect 2038 6332 2044 6384
rect 2096 6372 2102 6384
rect 2149 6375 2207 6381
rect 2149 6372 2161 6375
rect 2096 6344 2161 6372
rect 2096 6332 2102 6344
rect 2149 6341 2161 6344
rect 2195 6372 2207 6375
rect 3237 6375 3295 6381
rect 3237 6372 3249 6375
rect 2195 6344 3249 6372
rect 2195 6341 2207 6344
rect 2149 6335 2207 6341
rect 3237 6341 3249 6344
rect 3283 6341 3295 6375
rect 3237 6335 3295 6341
rect 3326 6332 3332 6384
rect 3384 6372 3390 6384
rect 4890 6372 4896 6384
rect 3384 6344 4896 6372
rect 3384 6332 3390 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 842 6060 848 6112
rect 900 6100 906 6112
rect 1489 6103 1547 6109
rect 1489 6100 1501 6103
rect 900 6072 1501 6100
rect 900 6060 906 6072
rect 1489 6069 1501 6072
rect 1535 6069 1547 6103
rect 1688 6100 1716 6267
rect 3418 6264 3424 6316
rect 3476 6264 3482 6316
rect 3528 6313 3556 6344
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 5074 6332 5080 6384
rect 5132 6381 5138 6384
rect 5132 6375 5151 6381
rect 5139 6341 5151 6375
rect 9950 6372 9956 6384
rect 5132 6335 5151 6341
rect 9600 6344 9956 6372
rect 5132 6332 5138 6335
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 3970 6304 3976 6316
rect 3927 6276 3976 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 9600 6313 9628 6344
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 10594 6332 10600 6384
rect 10652 6332 10658 6384
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 11422 6264 11428 6316
rect 11480 6304 11486 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 11480 6276 11529 6304
rect 11480 6264 11486 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 2590 6196 2596 6248
rect 2648 6236 2654 6248
rect 2685 6239 2743 6245
rect 2685 6236 2697 6239
rect 2648 6208 2697 6236
rect 2648 6196 2654 6208
rect 2685 6205 2697 6208
rect 2731 6205 2743 6239
rect 2685 6199 2743 6205
rect 2958 6168 2964 6180
rect 2148 6140 2964 6168
rect 2148 6109 2176 6140
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 3050 6128 3056 6180
rect 3108 6128 3114 6180
rect 3436 6168 3464 6264
rect 9398 6196 9404 6248
rect 9456 6196 9462 6248
rect 3436 6140 5120 6168
rect 2133 6103 2191 6109
rect 2133 6100 2145 6103
rect 1688 6072 2145 6100
rect 1489 6063 1547 6069
rect 2133 6069 2145 6072
rect 2179 6069 2191 6103
rect 2133 6063 2191 6069
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2590 6100 2596 6112
rect 2363 6072 2596 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 3142 6060 3148 6112
rect 3200 6060 3206 6112
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 3789 6103 3847 6109
rect 3789 6100 3801 6103
rect 3476 6072 3801 6100
rect 3476 6060 3482 6072
rect 3789 6069 3801 6072
rect 3835 6069 3847 6103
rect 3789 6063 3847 6069
rect 4065 6103 4123 6109
rect 4065 6069 4077 6103
rect 4111 6100 4123 6103
rect 4154 6100 4160 6112
rect 4111 6072 4160 6100
rect 4111 6069 4123 6072
rect 4065 6063 4123 6069
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 5092 6109 5120 6140
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 11204 6140 11744 6168
rect 11204 6128 11210 6140
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6069 5135 6103
rect 5077 6063 5135 6069
rect 5261 6103 5319 6109
rect 5261 6069 5273 6103
rect 5307 6100 5319 6103
rect 5350 6100 5356 6112
rect 5307 6072 5356 6100
rect 5307 6069 5319 6072
rect 5261 6063 5319 6069
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 9848 6103 9906 6109
rect 9848 6069 9860 6103
rect 9894 6100 9906 6103
rect 10042 6100 10048 6112
rect 9894 6072 10048 6100
rect 9894 6069 9906 6072
rect 9848 6063 9906 6069
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 11716 6109 11744 6140
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 11296 6072 11345 6100
rect 11296 6060 11302 6072
rect 11333 6069 11345 6072
rect 11379 6069 11391 6103
rect 11333 6063 11391 6069
rect 11701 6103 11759 6109
rect 11701 6069 11713 6103
rect 11747 6100 11759 6103
rect 12158 6100 12164 6112
rect 11747 6072 12164 6100
rect 11747 6069 11759 6072
rect 11701 6063 11759 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 1104 6010 12236 6032
rect 1104 5958 1550 6010
rect 1602 5958 1614 6010
rect 1666 5958 1678 6010
rect 1730 5958 1742 6010
rect 1794 5958 1806 6010
rect 1858 5958 3550 6010
rect 3602 5958 3614 6010
rect 3666 5958 3678 6010
rect 3730 5958 3742 6010
rect 3794 5958 3806 6010
rect 3858 5958 5550 6010
rect 5602 5958 5614 6010
rect 5666 5958 5678 6010
rect 5730 5958 5742 6010
rect 5794 5958 5806 6010
rect 5858 5958 7550 6010
rect 7602 5958 7614 6010
rect 7666 5958 7678 6010
rect 7730 5958 7742 6010
rect 7794 5958 7806 6010
rect 7858 5958 9550 6010
rect 9602 5958 9614 6010
rect 9666 5958 9678 6010
rect 9730 5958 9742 6010
rect 9794 5958 9806 6010
rect 9858 5958 11550 6010
rect 11602 5958 11614 6010
rect 11666 5958 11678 6010
rect 11730 5958 11742 6010
rect 11794 5958 11806 6010
rect 11858 5958 12236 6010
rect 1104 5936 12236 5958
rect 1946 5856 1952 5908
rect 2004 5856 2010 5908
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3605 5899 3663 5905
rect 3605 5896 3617 5899
rect 2924 5868 3617 5896
rect 2924 5856 2930 5868
rect 3605 5865 3617 5868
rect 3651 5865 3663 5899
rect 3605 5859 3663 5865
rect 9953 5899 10011 5905
rect 9953 5865 9965 5899
rect 9999 5896 10011 5899
rect 10042 5896 10048 5908
rect 9999 5868 10048 5896
rect 9999 5865 10011 5868
rect 9953 5859 10011 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 1964 5760 1992 5856
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 11609 5831 11667 5837
rect 11609 5828 11621 5831
rect 9824 5800 11621 5828
rect 9824 5788 9830 5800
rect 11609 5797 11621 5800
rect 11655 5797 11667 5831
rect 11609 5791 11667 5797
rect 2866 5760 2872 5772
rect 1688 5732 2872 5760
rect 1688 5701 1716 5732
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 3142 5720 3148 5772
rect 3200 5760 3206 5772
rect 5261 5763 5319 5769
rect 5261 5760 5273 5763
rect 3200 5732 5273 5760
rect 3200 5720 3206 5732
rect 5261 5729 5273 5732
rect 5307 5729 5319 5763
rect 8570 5760 8576 5772
rect 5261 5723 5319 5729
rect 8404 5732 8576 5760
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 842 5516 848 5568
rect 900 5556 906 5568
rect 1489 5559 1547 5565
rect 1489 5556 1501 5559
rect 900 5528 1501 5556
rect 900 5516 906 5528
rect 1489 5525 1501 5528
rect 1535 5525 1547 5559
rect 1872 5556 1900 5655
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5692 5595 5695
rect 5629 5695 5687 5701
rect 5629 5692 5641 5695
rect 5583 5664 5641 5692
rect 5583 5661 5595 5664
rect 5537 5655 5595 5661
rect 5629 5661 5641 5664
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 2130 5584 2136 5636
rect 2188 5584 2194 5636
rect 3418 5624 3424 5636
rect 3358 5596 3424 5624
rect 3418 5584 3424 5596
rect 3476 5584 3482 5636
rect 5552 5624 5580 5655
rect 7282 5652 7288 5704
rect 7340 5692 7346 5704
rect 8404 5701 8432 5732
rect 8570 5720 8576 5732
rect 8628 5760 8634 5772
rect 9030 5760 9036 5772
rect 8628 5732 9036 5760
rect 8628 5720 8634 5732
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10686 5760 10692 5772
rect 10459 5732 10692 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 10778 5720 10784 5772
rect 10836 5760 10842 5772
rect 10836 5732 11008 5760
rect 10836 5720 10842 5732
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 7340 5664 8033 5692
rect 7340 5652 7346 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 10321 5695 10379 5701
rect 8803 5664 10272 5692
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 5460 5596 5580 5624
rect 5460 5568 5488 5596
rect 5902 5584 5908 5636
rect 5960 5584 5966 5636
rect 7130 5596 7604 5624
rect 1946 5556 1952 5568
rect 1872 5528 1952 5556
rect 1489 5519 1547 5525
rect 1946 5516 1952 5528
rect 2004 5516 2010 5568
rect 2958 5516 2964 5568
rect 3016 5556 3022 5568
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 3016 5528 3801 5556
rect 3016 5516 3022 5528
rect 3789 5525 3801 5528
rect 3835 5556 3847 5559
rect 3878 5556 3884 5568
rect 3835 5528 3884 5556
rect 3835 5525 3847 5528
rect 3789 5519 3847 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 5442 5516 5448 5568
rect 5500 5516 5506 5568
rect 7282 5516 7288 5568
rect 7340 5556 7346 5568
rect 7377 5559 7435 5565
rect 7377 5556 7389 5559
rect 7340 5528 7389 5556
rect 7340 5516 7346 5528
rect 7377 5525 7389 5528
rect 7423 5525 7435 5559
rect 7377 5519 7435 5525
rect 7466 5516 7472 5568
rect 7524 5516 7530 5568
rect 7576 5556 7604 5596
rect 8110 5584 8116 5636
rect 8168 5624 8174 5636
rect 8941 5627 8999 5633
rect 8941 5624 8953 5627
rect 8168 5596 8953 5624
rect 8168 5584 8174 5596
rect 8941 5593 8953 5596
rect 8987 5624 8999 5627
rect 9950 5624 9956 5636
rect 8987 5596 9956 5624
rect 8987 5593 8999 5596
rect 8941 5587 8999 5593
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 10244 5624 10272 5664
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10873 5695 10931 5701
rect 10873 5692 10885 5695
rect 10367 5664 10885 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10873 5661 10885 5664
rect 10919 5661 10931 5695
rect 10980 5692 11008 5732
rect 11238 5720 11244 5772
rect 11296 5760 11302 5772
rect 11425 5763 11483 5769
rect 11425 5760 11437 5763
rect 11296 5732 11437 5760
rect 11296 5720 11302 5732
rect 11425 5729 11437 5732
rect 11471 5729 11483 5763
rect 11425 5723 11483 5729
rect 11885 5695 11943 5701
rect 11885 5692 11897 5695
rect 10980 5664 11897 5692
rect 10873 5655 10931 5661
rect 11885 5661 11897 5664
rect 11931 5661 11943 5695
rect 11885 5655 11943 5661
rect 10962 5624 10968 5636
rect 10244 5596 10968 5624
rect 10962 5584 10968 5596
rect 11020 5584 11026 5636
rect 11330 5584 11336 5636
rect 11388 5624 11394 5636
rect 11609 5627 11667 5633
rect 11609 5624 11621 5627
rect 11388 5596 11621 5624
rect 11388 5584 11394 5596
rect 11609 5593 11621 5596
rect 11655 5593 11667 5627
rect 11609 5587 11667 5593
rect 8297 5559 8355 5565
rect 8297 5556 8309 5559
rect 7576 5528 8309 5556
rect 8297 5525 8309 5528
rect 8343 5525 8355 5559
rect 8297 5519 8355 5525
rect 8662 5516 8668 5568
rect 8720 5516 8726 5568
rect 11790 5516 11796 5568
rect 11848 5516 11854 5568
rect 1104 5466 12236 5488
rect 1104 5414 2250 5466
rect 2302 5414 2314 5466
rect 2366 5414 2378 5466
rect 2430 5414 2442 5466
rect 2494 5414 2506 5466
rect 2558 5414 4250 5466
rect 4302 5414 4314 5466
rect 4366 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 6250 5466
rect 6302 5414 6314 5466
rect 6366 5414 6378 5466
rect 6430 5414 6442 5466
rect 6494 5414 6506 5466
rect 6558 5414 8250 5466
rect 8302 5414 8314 5466
rect 8366 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 10250 5466
rect 10302 5414 10314 5466
rect 10366 5414 10378 5466
rect 10430 5414 10442 5466
rect 10494 5414 10506 5466
rect 10558 5414 12236 5466
rect 1104 5392 12236 5414
rect 3878 5312 3884 5364
rect 3936 5312 3942 5364
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 4062 5352 4068 5364
rect 4019 5324 4068 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 5074 5352 5080 5364
rect 4295 5324 5080 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 5074 5312 5080 5324
rect 5132 5352 5138 5364
rect 5537 5355 5595 5361
rect 5537 5352 5549 5355
rect 5132 5324 5549 5352
rect 5132 5312 5138 5324
rect 5537 5321 5549 5324
rect 5583 5321 5595 5355
rect 5537 5315 5595 5321
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 5960 5324 6377 5352
rect 5960 5312 5966 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 9490 5312 9496 5364
rect 9548 5352 9554 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 9548 5324 9689 5352
rect 9548 5312 9554 5324
rect 9677 5321 9689 5324
rect 9723 5321 9735 5355
rect 9677 5315 9735 5321
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10134 5352 10140 5364
rect 9907 5324 10140 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 3326 5244 3332 5296
rect 3384 5284 3390 5296
rect 5445 5287 5503 5293
rect 5445 5284 5457 5287
rect 3384 5256 5457 5284
rect 3384 5244 3390 5256
rect 5445 5253 5457 5256
rect 5491 5253 5503 5287
rect 5445 5247 5503 5253
rect 5813 5287 5871 5293
rect 5813 5253 5825 5287
rect 5859 5284 5871 5287
rect 6914 5284 6920 5296
rect 5859 5256 6920 5284
rect 5859 5253 5871 5256
rect 5813 5247 5871 5253
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 1719 5188 2697 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 3237 5219 3295 5225
rect 3237 5216 3249 5219
rect 2924 5188 3249 5216
rect 2924 5176 2930 5188
rect 3237 5185 3249 5188
rect 3283 5216 3295 5219
rect 3418 5216 3424 5228
rect 3283 5188 3424 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 3418 5176 3424 5188
rect 3476 5216 3482 5228
rect 3697 5219 3755 5225
rect 3697 5216 3709 5219
rect 3476 5188 3709 5216
rect 3476 5176 3482 5188
rect 3697 5185 3709 5188
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 4614 5216 4620 5228
rect 4111 5188 4620 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4890 5176 4896 5228
rect 4948 5216 4954 5228
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 4948 5188 5273 5216
rect 4948 5176 4954 5188
rect 5261 5185 5273 5188
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 5902 5216 5908 5228
rect 5675 5188 5908 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 6564 5225 6592 5256
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 7466 5284 7472 5296
rect 7024 5256 7472 5284
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6822 5176 6828 5228
rect 6880 5176 6886 5228
rect 7024 5225 7052 5256
rect 7466 5244 7472 5256
rect 7524 5244 7530 5296
rect 8110 5284 8116 5296
rect 7944 5256 8116 5284
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 7944 5225 7972 5256
rect 8110 5244 8116 5256
rect 8168 5244 8174 5296
rect 8662 5244 8668 5296
rect 8720 5244 8726 5296
rect 9692 5284 9720 5315
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10413 5355 10471 5361
rect 10413 5321 10425 5355
rect 10459 5352 10471 5355
rect 10594 5352 10600 5364
rect 10459 5324 10600 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 10704 5324 11008 5352
rect 10704 5284 10732 5324
rect 10778 5293 10784 5296
rect 9692 5256 10732 5284
rect 10765 5287 10784 5293
rect 10765 5253 10777 5287
rect 10765 5247 10784 5253
rect 10778 5244 10784 5247
rect 10836 5244 10842 5296
rect 10980 5293 11008 5324
rect 11238 5312 11244 5364
rect 11296 5352 11302 5364
rect 11675 5355 11733 5361
rect 11675 5352 11687 5355
rect 11296 5324 11687 5352
rect 11296 5312 11302 5324
rect 11675 5321 11687 5324
rect 11721 5321 11733 5355
rect 11675 5315 11733 5321
rect 10965 5287 11023 5293
rect 10965 5253 10977 5287
rect 11011 5284 11023 5287
rect 11146 5284 11152 5296
rect 11011 5256 11152 5284
rect 11011 5253 11023 5256
rect 10965 5247 11023 5253
rect 11146 5244 11152 5256
rect 11204 5284 11210 5296
rect 11790 5284 11796 5296
rect 11204 5256 11796 5284
rect 11204 5244 11210 5256
rect 11790 5244 11796 5256
rect 11848 5284 11854 5296
rect 11885 5287 11943 5293
rect 11885 5284 11897 5287
rect 11848 5256 11897 5284
rect 11848 5244 11854 5256
rect 11885 5253 11897 5256
rect 11931 5253 11943 5287
rect 11885 5247 11943 5253
rect 7929 5219 7987 5225
rect 7929 5216 7941 5219
rect 7156 5188 7941 5216
rect 7156 5176 7162 5188
rect 7929 5185 7941 5188
rect 7975 5185 7987 5219
rect 7929 5179 7987 5185
rect 9766 5176 9772 5228
rect 9824 5176 9830 5228
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10134 5216 10140 5228
rect 10091 5188 10140 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5148 1823 5151
rect 1854 5148 1860 5160
rect 1811 5120 1860 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5148 2099 5151
rect 2130 5148 2136 5160
rect 2087 5120 2136 5148
rect 2087 5117 2099 5120
rect 2041 5111 2099 5117
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8938 5148 8944 5160
rect 8251 5120 8944 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8938 5108 8944 5120
rect 8996 5108 9002 5160
rect 9968 5148 9996 5179
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5216 10379 5219
rect 11054 5216 11060 5228
rect 10367 5188 11060 5216
rect 10367 5185 10379 5188
rect 10321 5179 10379 5185
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 12158 5216 12164 5228
rect 11379 5188 12164 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 9968 5120 10640 5148
rect 10612 5089 10640 5120
rect 10597 5083 10655 5089
rect 10597 5049 10609 5083
rect 10643 5080 10655 5083
rect 10686 5080 10692 5092
rect 10643 5052 10692 5080
rect 10643 5049 10655 5052
rect 10597 5043 10655 5049
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 11974 5080 11980 5092
rect 10796 5052 11980 5080
rect 10042 4972 10048 5024
rect 10100 5012 10106 5024
rect 10796 5021 10824 5052
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 10100 4984 10241 5012
rect 10100 4972 10106 4984
rect 10229 4981 10241 4984
rect 10275 4981 10287 5015
rect 10229 4975 10287 4981
rect 10781 5015 10839 5021
rect 10781 4981 10793 5015
rect 10827 4981 10839 5015
rect 10781 4975 10839 4981
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 11112 4984 11161 5012
rect 11112 4972 11118 4984
rect 11149 4981 11161 4984
rect 11195 4981 11207 5015
rect 11149 4975 11207 4981
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 11716 5021 11744 5052
rect 11974 5040 11980 5052
rect 12032 5040 12038 5092
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11388 4984 11529 5012
rect 11388 4972 11394 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 11701 5015 11759 5021
rect 11701 4981 11713 5015
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 1104 4922 12236 4944
rect 1104 4870 1550 4922
rect 1602 4870 1614 4922
rect 1666 4870 1678 4922
rect 1730 4870 1742 4922
rect 1794 4870 1806 4922
rect 1858 4870 3550 4922
rect 3602 4870 3614 4922
rect 3666 4870 3678 4922
rect 3730 4870 3742 4922
rect 3794 4870 3806 4922
rect 3858 4870 5550 4922
rect 5602 4870 5614 4922
rect 5666 4870 5678 4922
rect 5730 4870 5742 4922
rect 5794 4870 5806 4922
rect 5858 4870 7550 4922
rect 7602 4870 7614 4922
rect 7666 4870 7678 4922
rect 7730 4870 7742 4922
rect 7794 4870 7806 4922
rect 7858 4870 9550 4922
rect 9602 4870 9614 4922
rect 9666 4870 9678 4922
rect 9730 4870 9742 4922
rect 9794 4870 9806 4922
rect 9858 4870 11550 4922
rect 11602 4870 11614 4922
rect 11666 4870 11678 4922
rect 11730 4870 11742 4922
rect 11794 4870 11806 4922
rect 11858 4870 12236 4922
rect 1104 4848 12236 4870
rect 3050 4768 3056 4820
rect 3108 4768 3114 4820
rect 7374 4808 7380 4820
rect 6288 4780 7380 4808
rect 3326 4740 3332 4752
rect 3252 4712 3332 4740
rect 3252 4681 3280 4712
rect 3326 4700 3332 4712
rect 3384 4700 3390 4752
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 3418 4632 3424 4684
rect 3476 4632 3482 4684
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 3878 4672 3884 4684
rect 3559 4644 3884 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 5994 4632 6000 4684
rect 6052 4672 6058 4684
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 6052 4644 6193 4672
rect 6052 4632 6058 4644
rect 6181 4641 6193 4644
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 3326 4564 3332 4616
rect 3384 4564 3390 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 2590 4496 2596 4548
rect 2648 4536 2654 4548
rect 3988 4536 4016 4567
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 6288 4613 6316 4780
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 10008 4780 10241 4808
rect 10008 4768 10014 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10229 4771 10287 4777
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 10965 4811 11023 4817
rect 10965 4808 10977 4811
rect 10836 4780 10977 4808
rect 10836 4768 10842 4780
rect 10965 4777 10977 4780
rect 11011 4777 11023 4811
rect 10965 4771 11023 4777
rect 11793 4811 11851 4817
rect 11793 4777 11805 4811
rect 11839 4808 11851 4811
rect 11882 4808 11888 4820
rect 11839 4780 11888 4808
rect 11839 4777 11851 4780
rect 11793 4771 11851 4777
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 9490 4700 9496 4752
rect 9548 4740 9554 4752
rect 10796 4740 10824 4768
rect 9548 4712 10824 4740
rect 11425 4743 11483 4749
rect 9548 4700 9554 4712
rect 11425 4709 11437 4743
rect 11471 4740 11483 4743
rect 12066 4740 12072 4752
rect 11471 4712 12072 4740
rect 11471 4709 11483 4712
rect 11425 4703 11483 4709
rect 12066 4700 12072 4712
rect 12124 4700 12130 4752
rect 6641 4675 6699 4681
rect 6641 4641 6653 4675
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 6733 4675 6791 4681
rect 6733 4641 6745 4675
rect 6779 4672 6791 4675
rect 7098 4672 7104 4684
rect 6779 4644 7104 4672
rect 6779 4641 6791 4644
rect 6733 4635 6791 4641
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4573 6331 4607
rect 6656 4604 6684 4635
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8481 4675 8539 4681
rect 8481 4672 8493 4675
rect 8076 4644 8493 4672
rect 8076 4632 8082 4644
rect 8481 4641 8493 4644
rect 8527 4641 8539 4675
rect 8481 4635 8539 4641
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11204 4644 11652 4672
rect 11204 4632 11210 4644
rect 6656 4576 6776 4604
rect 6273 4567 6331 4573
rect 2648 4508 4016 4536
rect 4249 4539 4307 4545
rect 2648 4496 2654 4508
rect 4249 4505 4261 4539
rect 4295 4505 4307 4539
rect 4249 4499 4307 4505
rect 5997 4539 6055 4545
rect 5997 4505 6009 4539
rect 6043 4536 6055 4539
rect 6638 4536 6644 4548
rect 6043 4508 6644 4536
rect 6043 4505 6055 4508
rect 5997 4499 6055 4505
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 3292 4440 3801 4468
rect 3292 4428 3298 4440
rect 3789 4437 3801 4440
rect 3835 4437 3847 4471
rect 3789 4431 3847 4437
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4264 4468 4292 4499
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 6748 4536 6776 4576
rect 8110 4564 8116 4616
rect 8168 4564 8174 4616
rect 11238 4564 11244 4616
rect 11296 4564 11302 4616
rect 11624 4613 11652 4644
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 7009 4539 7067 4545
rect 7009 4536 7021 4539
rect 6748 4508 7021 4536
rect 7009 4505 7021 4508
rect 7055 4505 7067 4539
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 7009 4499 7067 4505
rect 8312 4508 8953 4536
rect 4212 4440 4292 4468
rect 6656 4468 6684 4496
rect 8312 4468 8340 4508
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 8941 4499 8999 4505
rect 9398 4496 9404 4548
rect 9456 4536 9462 4548
rect 9456 4508 10916 4536
rect 9456 4496 9462 4508
rect 6656 4440 8340 4468
rect 4212 4428 4218 4440
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10686 4468 10692 4480
rect 10284 4440 10692 4468
rect 10284 4428 10290 4440
rect 10686 4428 10692 4440
rect 10744 4468 10750 4480
rect 10781 4471 10839 4477
rect 10781 4468 10793 4471
rect 10744 4440 10793 4468
rect 10744 4428 10750 4440
rect 10781 4437 10793 4440
rect 10827 4437 10839 4471
rect 10888 4468 10916 4508
rect 11146 4496 11152 4548
rect 11204 4496 11210 4548
rect 10949 4471 11007 4477
rect 10949 4468 10961 4471
rect 10888 4440 10961 4468
rect 10781 4431 10839 4437
rect 10949 4437 10961 4440
rect 10995 4468 11007 4471
rect 11330 4468 11336 4480
rect 10995 4440 11336 4468
rect 10995 4437 11007 4440
rect 10949 4431 11007 4437
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 1104 4378 12236 4400
rect 1104 4326 2250 4378
rect 2302 4326 2314 4378
rect 2366 4326 2378 4378
rect 2430 4326 2442 4378
rect 2494 4326 2506 4378
rect 2558 4326 4250 4378
rect 4302 4326 4314 4378
rect 4366 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 6250 4378
rect 6302 4326 6314 4378
rect 6366 4326 6378 4378
rect 6430 4326 6442 4378
rect 6494 4326 6506 4378
rect 6558 4326 8250 4378
rect 8302 4326 8314 4378
rect 8366 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 10250 4378
rect 10302 4326 10314 4378
rect 10366 4326 10378 4378
rect 10430 4326 10442 4378
rect 10494 4326 10506 4378
rect 10558 4326 12236 4378
rect 1104 4304 12236 4326
rect 5629 4267 5687 4273
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 5718 4264 5724 4276
rect 5675 4236 5724 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 5813 4267 5871 4273
rect 5813 4233 5825 4267
rect 5859 4264 5871 4267
rect 7282 4264 7288 4276
rect 5859 4236 7288 4264
rect 5859 4233 5871 4236
rect 5813 4227 5871 4233
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 9398 4264 9404 4276
rect 8864 4236 9404 4264
rect 5997 4199 6055 4205
rect 5997 4165 6009 4199
rect 6043 4196 6055 4199
rect 6086 4196 6092 4208
rect 6043 4168 6092 4196
rect 6043 4165 6055 4168
rect 5997 4159 6055 4165
rect 6086 4156 6092 4168
rect 6144 4156 6150 4208
rect 6914 4196 6920 4208
rect 6196 4168 6920 4196
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 3513 4131 3571 4137
rect 3513 4128 3525 4131
rect 2363 4100 3525 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 3513 4097 3525 4100
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4212 4100 4261 4128
rect 4212 4088 4218 4100
rect 4249 4097 4261 4100
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 6196 4128 6224 4168
rect 6914 4156 6920 4168
rect 6972 4196 6978 4208
rect 6972 4168 8064 4196
rect 6972 4156 6978 4168
rect 8036 4140 8064 4168
rect 5951 4126 6040 4128
rect 6104 4126 6224 4128
rect 5951 4100 6224 4126
rect 6840 4100 7052 4128
rect 5951 4097 5963 4100
rect 6012 4098 6132 4100
rect 5905 4091 5963 4097
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 3234 4060 3240 4072
rect 2455 4032 3240 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 3970 4060 3976 4072
rect 3476 4032 3976 4060
rect 3476 4020 3482 4032
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4060 4123 4063
rect 4614 4060 4620 4072
rect 4111 4032 4620 4060
rect 4111 4029 4123 4032
rect 4065 4023 4123 4029
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 5552 4060 5580 4091
rect 6840 4060 6868 4100
rect 5552 4032 6868 4060
rect 6917 4063 6975 4069
rect 3878 3952 3884 4004
rect 3936 3992 3942 4004
rect 4246 3992 4252 4004
rect 3936 3964 4252 3992
rect 3936 3952 3942 3964
rect 4246 3952 4252 3964
rect 4304 3992 4310 4004
rect 5552 3992 5580 4032
rect 6917 4029 6929 4063
rect 6963 4029 6975 4063
rect 7024 4060 7052 4100
rect 7374 4088 7380 4140
rect 7432 4088 7438 4140
rect 8018 4088 8024 4140
rect 8076 4088 8082 4140
rect 8864 4137 8892 4236
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 9490 4224 9496 4276
rect 9548 4224 9554 4276
rect 9585 4267 9643 4273
rect 9585 4233 9597 4267
rect 9631 4264 9643 4267
rect 10410 4264 10416 4276
rect 9631 4236 10416 4264
rect 9631 4233 9643 4236
rect 9585 4227 9643 4233
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 9125 4199 9183 4205
rect 9125 4165 9137 4199
rect 9171 4196 9183 4199
rect 10597 4199 10655 4205
rect 10597 4196 10609 4199
rect 9171 4168 10609 4196
rect 9171 4165 9183 4168
rect 9125 4159 9183 4165
rect 10597 4165 10609 4168
rect 10643 4165 10655 4199
rect 10597 4159 10655 4165
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 9490 4128 9496 4140
rect 8987 4100 9496 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 7024 4032 8401 4060
rect 6917 4023 6975 4029
rect 8389 4029 8401 4032
rect 8435 4060 8447 4063
rect 8478 4060 8484 4072
rect 8435 4032 8484 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 4304 3964 5580 3992
rect 4304 3952 4310 3964
rect 6178 3952 6184 4004
rect 6236 3992 6242 4004
rect 6932 3992 6960 4023
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 6236 3964 6960 3992
rect 8588 3992 8616 4091
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4128 9827 4131
rect 11146 4128 11152 4140
rect 9815 4100 11152 4128
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 11146 4088 11152 4100
rect 11204 4128 11210 4140
rect 11609 4131 11667 4137
rect 11609 4128 11621 4131
rect 11204 4100 11621 4128
rect 11204 4088 11210 4100
rect 11609 4097 11621 4100
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 9052 4063 9110 4069
rect 9052 4029 9064 4063
rect 9098 4060 9110 4063
rect 10134 4060 10140 4072
rect 9098 4032 10140 4060
rect 9098 4029 9110 4032
rect 9052 4023 9110 4029
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 10410 4020 10416 4072
rect 10468 4020 10474 4072
rect 12158 4060 12164 4072
rect 11716 4032 12164 4060
rect 11716 3992 11744 4032
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 8588 3964 11744 3992
rect 6236 3952 6242 3964
rect 11790 3952 11796 4004
rect 11848 3952 11854 4004
rect 2682 3884 2688 3936
rect 2740 3884 2746 3936
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 5166 3884 5172 3936
rect 5224 3924 5230 3936
rect 5445 3927 5503 3933
rect 5445 3924 5457 3927
rect 5224 3896 5457 3924
rect 5224 3884 5230 3896
rect 5445 3893 5457 3896
rect 5491 3893 5503 3927
rect 5445 3887 5503 3893
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 5960 3896 6377 3924
rect 5960 3884 5966 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 9214 3884 9220 3936
rect 9272 3884 9278 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9456 3896 9873 3924
rect 9456 3884 9462 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 1104 3834 12236 3856
rect 1104 3782 1550 3834
rect 1602 3782 1614 3834
rect 1666 3782 1678 3834
rect 1730 3782 1742 3834
rect 1794 3782 1806 3834
rect 1858 3782 3550 3834
rect 3602 3782 3614 3834
rect 3666 3782 3678 3834
rect 3730 3782 3742 3834
rect 3794 3782 3806 3834
rect 3858 3782 5550 3834
rect 5602 3782 5614 3834
rect 5666 3782 5678 3834
rect 5730 3782 5742 3834
rect 5794 3782 5806 3834
rect 5858 3782 7550 3834
rect 7602 3782 7614 3834
rect 7666 3782 7678 3834
rect 7730 3782 7742 3834
rect 7794 3782 7806 3834
rect 7858 3782 9550 3834
rect 9602 3782 9614 3834
rect 9666 3782 9678 3834
rect 9730 3782 9742 3834
rect 9794 3782 9806 3834
rect 9858 3782 11550 3834
rect 11602 3782 11614 3834
rect 11666 3782 11678 3834
rect 11730 3782 11742 3834
rect 11794 3782 11806 3834
rect 11858 3782 12236 3834
rect 1104 3760 12236 3782
rect 1946 3680 1952 3732
rect 2004 3680 2010 3732
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 6052 3692 7849 3720
rect 6052 3680 6058 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 7837 3683 7895 3689
rect 8021 3723 8079 3729
rect 8021 3689 8033 3723
rect 8067 3689 8079 3723
rect 8021 3683 8079 3689
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 1964 3584 1992 3680
rect 8036 3652 8064 3683
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 8168 3692 8493 3720
rect 8168 3680 8174 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 10686 3720 10692 3732
rect 8481 3683 8539 3689
rect 9324 3692 10692 3720
rect 7760 3624 8064 3652
rect 4154 3584 4160 3596
rect 1903 3556 4160 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 4154 3544 4160 3556
rect 4212 3584 4218 3596
rect 5442 3584 5448 3596
rect 4212 3556 5448 3584
rect 4212 3544 4218 3556
rect 5442 3544 5448 3556
rect 5500 3584 5506 3596
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 5500 3556 6009 3584
rect 5500 3544 5506 3556
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 6270 3544 6276 3596
rect 6328 3584 6334 3596
rect 6730 3584 6736 3596
rect 6328 3556 6736 3584
rect 6328 3544 6334 3556
rect 6730 3544 6736 3556
rect 6788 3584 6794 3596
rect 7760 3593 7788 3624
rect 9324 3593 9352 3692
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 11425 3723 11483 3729
rect 11425 3720 11437 3723
rect 11204 3692 11437 3720
rect 11204 3680 11210 3692
rect 11425 3689 11437 3692
rect 11471 3689 11483 3723
rect 11425 3683 11483 3689
rect 7745 3587 7803 3593
rect 7745 3584 7757 3587
rect 6788 3556 7757 3584
rect 6788 3544 6794 3556
rect 7745 3553 7757 3556
rect 7791 3553 7803 3587
rect 7745 3547 7803 3553
rect 9309 3587 9367 3593
rect 9309 3553 9321 3587
rect 9355 3553 9367 3587
rect 9309 3547 9367 3553
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 9950 3584 9956 3596
rect 9723 3556 9956 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 2130 3408 2136 3460
rect 2188 3408 2194 3460
rect 3881 3451 3939 3457
rect 3881 3448 3893 3451
rect 3358 3420 3893 3448
rect 3881 3417 3893 3420
rect 3927 3417 3939 3451
rect 3988 3448 4016 3479
rect 7374 3476 7380 3528
rect 7432 3476 7438 3528
rect 8018 3476 8024 3528
rect 8076 3516 8082 3528
rect 8478 3516 8484 3528
rect 8076 3488 8484 3516
rect 8076 3476 8082 3488
rect 8478 3476 8484 3488
rect 8536 3516 8542 3528
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 8536 3488 8585 3516
rect 8536 3476 8542 3488
rect 8573 3485 8585 3488
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9398 3516 9404 3528
rect 9263 3488 9404 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 4154 3448 4160 3460
rect 3988 3420 4160 3448
rect 3881 3411 3939 3417
rect 4154 3408 4160 3420
rect 4212 3408 4218 3460
rect 4433 3451 4491 3457
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 4706 3448 4712 3460
rect 4479 3420 4712 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 5166 3408 5172 3460
rect 5224 3408 5230 3460
rect 6178 3448 6184 3460
rect 5920 3420 6184 3448
rect 3418 3340 3424 3392
rect 3476 3380 3482 3392
rect 3605 3383 3663 3389
rect 3605 3380 3617 3383
rect 3476 3352 3617 3380
rect 3476 3340 3482 3352
rect 3605 3349 3617 3352
rect 3651 3349 3663 3383
rect 3605 3343 3663 3349
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 5920 3389 5948 3420
rect 6178 3408 6184 3420
rect 6236 3408 6242 3460
rect 6273 3451 6331 3457
rect 6273 3417 6285 3451
rect 6319 3417 6331 3451
rect 8205 3451 8263 3457
rect 8205 3448 8217 3451
rect 6273 3411 6331 3417
rect 7576 3420 8217 3448
rect 5905 3383 5963 3389
rect 5905 3380 5917 3383
rect 5868 3352 5917 3380
rect 5868 3340 5874 3352
rect 5905 3349 5917 3352
rect 5951 3349 5963 3383
rect 5905 3343 5963 3349
rect 6086 3340 6092 3392
rect 6144 3380 6150 3392
rect 6288 3380 6316 3411
rect 6144 3352 6316 3380
rect 6144 3340 6150 3352
rect 6362 3340 6368 3392
rect 6420 3380 6426 3392
rect 7576 3380 7604 3420
rect 8205 3417 8217 3420
rect 8251 3417 8263 3451
rect 9600 3448 9628 3547
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10410 3544 10416 3596
rect 10468 3584 10474 3596
rect 10962 3584 10968 3596
rect 10468 3556 10968 3584
rect 10468 3544 10474 3556
rect 10962 3544 10968 3556
rect 11020 3584 11026 3596
rect 11020 3556 11652 3584
rect 11020 3544 11026 3556
rect 11624 3525 11652 3556
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 9858 3448 9864 3460
rect 9600 3420 9864 3448
rect 8205 3411 8263 3417
rect 9858 3408 9864 3420
rect 9916 3408 9922 3460
rect 9953 3451 10011 3457
rect 9953 3417 9965 3451
rect 9999 3448 10011 3451
rect 10042 3448 10048 3460
rect 9999 3420 10048 3448
rect 9999 3417 10011 3420
rect 9953 3411 10011 3417
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 10686 3408 10692 3460
rect 10744 3408 10750 3460
rect 6420 3352 7604 3380
rect 6420 3340 6426 3352
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 7995 3383 8053 3389
rect 7995 3380 8007 3383
rect 7708 3352 8007 3380
rect 7708 3340 7714 3352
rect 7995 3349 8007 3352
rect 8041 3349 8053 3383
rect 7995 3343 8053 3349
rect 11790 3340 11796 3392
rect 11848 3340 11854 3392
rect 1104 3290 12236 3312
rect 1104 3238 2250 3290
rect 2302 3238 2314 3290
rect 2366 3238 2378 3290
rect 2430 3238 2442 3290
rect 2494 3238 2506 3290
rect 2558 3238 4250 3290
rect 4302 3238 4314 3290
rect 4366 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 6250 3290
rect 6302 3238 6314 3290
rect 6366 3238 6378 3290
rect 6430 3238 6442 3290
rect 6494 3238 6506 3290
rect 6558 3238 8250 3290
rect 8302 3238 8314 3290
rect 8366 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 10250 3290
rect 10302 3238 10314 3290
rect 10366 3238 10378 3290
rect 10430 3238 10442 3290
rect 10494 3238 10506 3290
rect 10558 3238 12236 3290
rect 1104 3216 12236 3238
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 2740 3148 3188 3176
rect 2740 3136 2746 3148
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 3160 3117 3188 3148
rect 4614 3136 4620 3188
rect 4672 3136 4678 3188
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 6733 3179 6791 3185
rect 5408 3148 6684 3176
rect 5408 3136 5414 3148
rect 3145 3111 3203 3117
rect 2004 3080 2912 3108
rect 2004 3068 2010 3080
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 2774 3040 2780 3052
rect 2363 3012 2780 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 2884 3049 2912 3080
rect 3145 3077 3157 3111
rect 3191 3077 3203 3111
rect 4430 3108 4436 3120
rect 4370 3080 4436 3108
rect 3145 3071 3203 3077
rect 4430 3068 4436 3080
rect 4488 3068 4494 3120
rect 5902 3108 5908 3120
rect 5276 3080 5908 3108
rect 5276 3049 5304 3080
rect 5902 3068 5908 3080
rect 5960 3068 5966 3120
rect 5994 3068 6000 3120
rect 6052 3108 6058 3120
rect 6656 3108 6684 3148
rect 6733 3145 6745 3179
rect 6779 3176 6791 3179
rect 6822 3176 6828 3188
rect 6779 3148 6828 3176
rect 6779 3145 6791 3148
rect 6733 3139 6791 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7668 3148 9628 3176
rect 7098 3108 7104 3120
rect 6052 3080 6592 3108
rect 6656 3080 7104 3108
rect 6052 3068 6058 3080
rect 6564 3049 6592 3080
rect 7098 3068 7104 3080
rect 7156 3108 7162 3120
rect 7558 3108 7564 3120
rect 7156 3080 7564 3108
rect 7156 3068 7162 3080
rect 7558 3068 7564 3080
rect 7616 3068 7622 3120
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3040 5779 3043
rect 6549 3043 6607 3049
rect 5767 3012 6500 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2130 2972 2136 2984
rect 1995 2944 2136 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 2590 2972 2596 2984
rect 2455 2944 2596 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 4706 2932 4712 2984
rect 4764 2972 4770 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4764 2944 4905 2972
rect 4764 2932 4770 2944
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 5350 2932 5356 2984
rect 5408 2932 5414 2984
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2941 5871 2975
rect 5813 2935 5871 2941
rect 5828 2904 5856 2935
rect 6362 2932 6368 2984
rect 6420 2932 6426 2984
rect 6472 2972 6500 3012
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 7668 3049 7696 3148
rect 9600 3108 9628 3148
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 11480 3148 11529 3176
rect 11480 3136 11486 3148
rect 11517 3145 11529 3148
rect 11563 3145 11575 3179
rect 11517 3139 11575 3145
rect 9950 3108 9956 3120
rect 9600 3080 9956 3108
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 6788 3012 7389 3040
rect 6788 3000 6794 3012
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9600 3049 9628 3080
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 11238 3108 11244 3120
rect 11086 3080 11244 3108
rect 11238 3068 11244 3080
rect 11296 3068 11302 3120
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3040 11759 3043
rect 11974 3040 11980 3052
rect 11747 3012 11980 3040
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6472 2944 6837 2972
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7926 2932 7932 2984
rect 7984 2932 7990 2984
rect 9858 2932 9864 2984
rect 9916 2932 9922 2984
rect 7006 2904 7012 2916
rect 5828 2876 7012 2904
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 11333 2907 11391 2913
rect 11333 2904 11345 2907
rect 11020 2876 11345 2904
rect 11020 2864 11026 2876
rect 11333 2873 11345 2876
rect 11379 2873 11391 2907
rect 11333 2867 11391 2873
rect 5997 2839 6055 2845
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 6086 2836 6092 2848
rect 6043 2808 6092 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6086 2796 6092 2808
rect 6144 2796 6150 2848
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 6914 2836 6920 2848
rect 6420 2808 6920 2836
rect 6420 2796 6426 2808
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 9950 2836 9956 2848
rect 9447 2808 9956 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 1104 2746 12236 2768
rect 1104 2694 1550 2746
rect 1602 2694 1614 2746
rect 1666 2694 1678 2746
rect 1730 2694 1742 2746
rect 1794 2694 1806 2746
rect 1858 2694 3550 2746
rect 3602 2694 3614 2746
rect 3666 2694 3678 2746
rect 3730 2694 3742 2746
rect 3794 2694 3806 2746
rect 3858 2694 5550 2746
rect 5602 2694 5614 2746
rect 5666 2694 5678 2746
rect 5730 2694 5742 2746
rect 5794 2694 5806 2746
rect 5858 2694 7550 2746
rect 7602 2694 7614 2746
rect 7666 2694 7678 2746
rect 7730 2694 7742 2746
rect 7794 2694 7806 2746
rect 7858 2694 9550 2746
rect 9602 2694 9614 2746
rect 9666 2694 9678 2746
rect 9730 2694 9742 2746
rect 9794 2694 9806 2746
rect 9858 2694 11550 2746
rect 11602 2694 11614 2746
rect 11666 2694 11678 2746
rect 11730 2694 11742 2746
rect 11794 2694 11806 2746
rect 11858 2694 12236 2746
rect 1104 2672 12236 2694
rect 4430 2592 4436 2644
rect 4488 2592 4494 2644
rect 7006 2592 7012 2644
rect 7064 2592 7070 2644
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 7653 2635 7711 2641
rect 7653 2632 7665 2635
rect 7432 2604 7665 2632
rect 7432 2592 7438 2604
rect 7653 2601 7665 2604
rect 7699 2601 7711 2635
rect 7653 2595 7711 2601
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8205 2635 8263 2641
rect 8205 2632 8217 2635
rect 7984 2604 8217 2632
rect 7984 2592 7990 2604
rect 8205 2601 8217 2604
rect 8251 2601 8263 2635
rect 8205 2595 8263 2601
rect 9030 2592 9036 2644
rect 9088 2592 9094 2644
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 10744 2604 10977 2632
rect 10744 2592 10750 2604
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 10965 2595 11023 2601
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 11974 2632 11980 2644
rect 11931 2604 11980 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 6914 2524 6920 2576
rect 6972 2564 6978 2576
rect 6972 2536 8156 2564
rect 6972 2524 6978 2536
rect 4614 2496 4620 2508
rect 4264 2468 4620 2496
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 4264 2437 4292 2468
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6052 2468 6960 2496
rect 6052 2456 6058 2468
rect 6196 2437 6224 2468
rect 3605 2431 3663 2437
rect 3605 2428 3617 2431
rect 3476 2400 3617 2428
rect 3476 2388 3482 2400
rect 3605 2397 3617 2400
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2428 6239 2431
rect 6227 2400 6261 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 4540 2360 4568 2391
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 6932 2437 6960 2468
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6788 2400 6837 2428
rect 6788 2388 6794 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7098 2388 7104 2440
rect 7156 2388 7162 2440
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7340 2400 7481 2428
rect 7340 2388 7346 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 8018 2428 8024 2440
rect 7791 2400 8024 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8128 2437 8156 2536
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 9214 2496 9220 2508
rect 8711 2468 9220 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 9950 2456 9956 2508
rect 10008 2456 10014 2508
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9968 2428 9996 2456
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9171 2400 9904 2428
rect 9968 2400 10149 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 4212 2332 4568 2360
rect 8588 2360 8616 2391
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8588 2332 9413 2360
rect 4212 2320 4218 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9876 2360 9904 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 11112 2400 11161 2428
rect 11112 2388 11118 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11072 2360 11100 2388
rect 9876 2332 11100 2360
rect 9401 2323 9459 2329
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3421 2295 3479 2301
rect 3421 2292 3433 2295
rect 3292 2264 3433 2292
rect 3292 2252 3298 2264
rect 3421 2261 3433 2264
rect 3467 2261 3479 2295
rect 3421 2255 3479 2261
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3936 2264 4077 2292
rect 3936 2252 3942 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 5997 2295 6055 2301
rect 5997 2292 6009 2295
rect 5868 2264 6009 2292
rect 5868 2252 5874 2264
rect 5997 2261 6009 2264
rect 6043 2261 6055 2295
rect 5997 2255 6055 2261
rect 6638 2252 6644 2304
rect 6696 2252 6702 2304
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 7156 2264 7297 2292
rect 7156 2252 7162 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7800 2264 7941 2292
rect 7800 2252 7806 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 10321 2295 10379 2301
rect 10321 2292 10333 2295
rect 9088 2264 10333 2292
rect 9088 2252 9094 2264
rect 10321 2261 10333 2264
rect 10367 2261 10379 2295
rect 10321 2255 10379 2261
rect 1104 2202 12236 2224
rect 1104 2150 2250 2202
rect 2302 2150 2314 2202
rect 2366 2150 2378 2202
rect 2430 2150 2442 2202
rect 2494 2150 2506 2202
rect 2558 2150 4250 2202
rect 4302 2150 4314 2202
rect 4366 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 6250 2202
rect 6302 2150 6314 2202
rect 6366 2150 6378 2202
rect 6430 2150 6442 2202
rect 6494 2150 6506 2202
rect 6558 2150 8250 2202
rect 8302 2150 8314 2202
rect 8366 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 10250 2202
rect 10302 2150 10314 2202
rect 10366 2150 10378 2202
rect 10430 2150 10442 2202
rect 10494 2150 10506 2202
rect 10558 2150 12236 2202
rect 1104 2128 12236 2150
<< via1 >>
rect 2250 13030 2302 13082
rect 2314 13030 2366 13082
rect 2378 13030 2430 13082
rect 2442 13030 2494 13082
rect 2506 13030 2558 13082
rect 4250 13030 4302 13082
rect 4314 13030 4366 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 6250 13030 6302 13082
rect 6314 13030 6366 13082
rect 6378 13030 6430 13082
rect 6442 13030 6494 13082
rect 6506 13030 6558 13082
rect 8250 13030 8302 13082
rect 8314 13030 8366 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 10250 13030 10302 13082
rect 10314 13030 10366 13082
rect 10378 13030 10430 13082
rect 10442 13030 10494 13082
rect 10506 13030 10558 13082
rect 4620 12928 4672 12980
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 6092 12971 6144 12980
rect 6092 12937 6101 12971
rect 6101 12937 6135 12971
rect 6135 12937 6144 12971
rect 6092 12928 6144 12937
rect 6736 12971 6788 12980
rect 6736 12937 6745 12971
rect 6745 12937 6779 12971
rect 6779 12937 6788 12971
rect 6736 12928 6788 12937
rect 11060 12860 11112 12912
rect 5264 12792 5316 12844
rect 5816 12792 5868 12844
rect 6000 12792 6052 12844
rect 6644 12792 6696 12844
rect 9956 12792 10008 12844
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 5172 12724 5224 12776
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 11244 12792 11296 12844
rect 12072 12792 12124 12844
rect 7380 12656 7432 12708
rect 10784 12656 10836 12708
rect 10140 12588 10192 12640
rect 11152 12588 11204 12640
rect 11336 12631 11388 12640
rect 11336 12597 11345 12631
rect 11345 12597 11379 12631
rect 11379 12597 11388 12631
rect 11336 12588 11388 12597
rect 11980 12588 12032 12640
rect 1550 12486 1602 12538
rect 1614 12486 1666 12538
rect 1678 12486 1730 12538
rect 1742 12486 1794 12538
rect 1806 12486 1858 12538
rect 3550 12486 3602 12538
rect 3614 12486 3666 12538
rect 3678 12486 3730 12538
rect 3742 12486 3794 12538
rect 3806 12486 3858 12538
rect 5550 12486 5602 12538
rect 5614 12486 5666 12538
rect 5678 12486 5730 12538
rect 5742 12486 5794 12538
rect 5806 12486 5858 12538
rect 7550 12486 7602 12538
rect 7614 12486 7666 12538
rect 7678 12486 7730 12538
rect 7742 12486 7794 12538
rect 7806 12486 7858 12538
rect 9550 12486 9602 12538
rect 9614 12486 9666 12538
rect 9678 12486 9730 12538
rect 9742 12486 9794 12538
rect 9806 12486 9858 12538
rect 11550 12486 11602 12538
rect 11614 12486 11666 12538
rect 11678 12486 11730 12538
rect 11742 12486 11794 12538
rect 11806 12486 11858 12538
rect 5448 12427 5500 12436
rect 5448 12393 5457 12427
rect 5457 12393 5491 12427
rect 5491 12393 5500 12427
rect 5448 12384 5500 12393
rect 5908 12427 5960 12436
rect 5908 12393 5917 12427
rect 5917 12393 5951 12427
rect 5951 12393 5960 12427
rect 5908 12384 5960 12393
rect 12072 12384 12124 12436
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 3884 12180 3936 12232
rect 5264 12180 5316 12232
rect 6644 12248 6696 12300
rect 10600 12316 10652 12368
rect 10048 12248 10100 12300
rect 6920 12180 6972 12232
rect 9312 12180 9364 12232
rect 9956 12180 10008 12232
rect 11428 12180 11480 12232
rect 10324 12112 10376 12164
rect 10692 12112 10744 12164
rect 4068 12087 4120 12096
rect 4068 12053 4077 12087
rect 4077 12053 4111 12087
rect 4111 12053 4120 12087
rect 4068 12044 4120 12053
rect 4160 12044 4212 12096
rect 5908 12044 5960 12096
rect 7196 12087 7248 12096
rect 7196 12053 7205 12087
rect 7205 12053 7239 12087
rect 7239 12053 7248 12087
rect 7196 12044 7248 12053
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 10048 12087 10100 12096
rect 10048 12053 10075 12087
rect 10075 12053 10100 12087
rect 10048 12044 10100 12053
rect 12164 12044 12216 12096
rect 2250 11942 2302 11994
rect 2314 11942 2366 11994
rect 2378 11942 2430 11994
rect 2442 11942 2494 11994
rect 2506 11942 2558 11994
rect 4250 11942 4302 11994
rect 4314 11942 4366 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 6250 11942 6302 11994
rect 6314 11942 6366 11994
rect 6378 11942 6430 11994
rect 6442 11942 6494 11994
rect 6506 11942 6558 11994
rect 8250 11942 8302 11994
rect 8314 11942 8366 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 10250 11942 10302 11994
rect 10314 11942 10366 11994
rect 10378 11942 10430 11994
rect 10442 11942 10494 11994
rect 10506 11942 10558 11994
rect 4160 11840 4212 11892
rect 5448 11840 5500 11892
rect 4068 11772 4120 11824
rect 3056 11679 3108 11688
rect 3056 11645 3065 11679
rect 3065 11645 3099 11679
rect 3099 11645 3108 11679
rect 3056 11636 3108 11645
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 7196 11772 7248 11824
rect 9496 11772 9548 11824
rect 10968 11772 11020 11824
rect 5908 11747 5960 11756
rect 5908 11713 5917 11747
rect 5917 11713 5951 11747
rect 5951 11713 5960 11747
rect 5908 11704 5960 11713
rect 10048 11704 10100 11756
rect 10876 11704 10928 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11336 11815 11388 11824
rect 11336 11781 11345 11815
rect 11345 11781 11379 11815
rect 11379 11781 11388 11815
rect 11336 11772 11388 11781
rect 6000 11636 6052 11688
rect 7380 11636 7432 11688
rect 5172 11568 5224 11620
rect 3976 11500 4028 11552
rect 5356 11500 5408 11552
rect 6644 11568 6696 11620
rect 6092 11543 6144 11552
rect 6092 11509 6101 11543
rect 6101 11509 6135 11543
rect 6135 11509 6144 11543
rect 6092 11500 6144 11509
rect 7104 11500 7156 11552
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 9220 11636 9272 11688
rect 10692 11636 10744 11688
rect 10048 11568 10100 11620
rect 11244 11568 11296 11620
rect 9956 11500 10008 11552
rect 11888 11500 11940 11552
rect 1550 11398 1602 11450
rect 1614 11398 1666 11450
rect 1678 11398 1730 11450
rect 1742 11398 1794 11450
rect 1806 11398 1858 11450
rect 3550 11398 3602 11450
rect 3614 11398 3666 11450
rect 3678 11398 3730 11450
rect 3742 11398 3794 11450
rect 3806 11398 3858 11450
rect 5550 11398 5602 11450
rect 5614 11398 5666 11450
rect 5678 11398 5730 11450
rect 5742 11398 5794 11450
rect 5806 11398 5858 11450
rect 7550 11398 7602 11450
rect 7614 11398 7666 11450
rect 7678 11398 7730 11450
rect 7742 11398 7794 11450
rect 7806 11398 7858 11450
rect 9550 11398 9602 11450
rect 9614 11398 9666 11450
rect 9678 11398 9730 11450
rect 9742 11398 9794 11450
rect 9806 11398 9858 11450
rect 11550 11398 11602 11450
rect 11614 11398 11666 11450
rect 11678 11398 11730 11450
rect 11742 11398 11794 11450
rect 11806 11398 11858 11450
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 5448 11296 5500 11348
rect 6920 11296 6972 11348
rect 8760 11296 8812 11348
rect 12072 11296 12124 11348
rect 3976 11203 4028 11212
rect 3976 11169 3985 11203
rect 3985 11169 4019 11203
rect 4019 11169 4028 11203
rect 3976 11160 4028 11169
rect 4620 11160 4672 11212
rect 5356 11228 5408 11280
rect 6000 11160 6052 11212
rect 6092 11160 6144 11212
rect 10140 11228 10192 11280
rect 5172 11092 5224 11144
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 8576 11160 8628 11212
rect 9220 11203 9272 11212
rect 9220 11169 9229 11203
rect 9229 11169 9263 11203
rect 9263 11169 9272 11203
rect 9220 11160 9272 11169
rect 10048 11160 10100 11212
rect 9956 11092 10008 11144
rect 5264 11024 5316 11076
rect 1952 10956 2004 11008
rect 3976 10956 4028 11008
rect 11060 11024 11112 11076
rect 2250 10854 2302 10906
rect 2314 10854 2366 10906
rect 2378 10854 2430 10906
rect 2442 10854 2494 10906
rect 2506 10854 2558 10906
rect 4250 10854 4302 10906
rect 4314 10854 4366 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 6250 10854 6302 10906
rect 6314 10854 6366 10906
rect 6378 10854 6430 10906
rect 6442 10854 6494 10906
rect 6506 10854 6558 10906
rect 8250 10854 8302 10906
rect 8314 10854 8366 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 10250 10854 10302 10906
rect 10314 10854 10366 10906
rect 10378 10854 10430 10906
rect 10442 10854 10494 10906
rect 10506 10854 10558 10906
rect 6000 10752 6052 10804
rect 11428 10752 11480 10804
rect 12164 10752 12216 10804
rect 3056 10684 3108 10736
rect 2688 10616 2740 10668
rect 4068 10684 4120 10736
rect 4896 10684 4948 10736
rect 8760 10616 8812 10668
rect 9036 10616 9088 10668
rect 9956 10684 10008 10736
rect 11152 10684 11204 10736
rect 4620 10548 4672 10600
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 10600 10548 10652 10600
rect 11060 10548 11112 10600
rect 848 10412 900 10464
rect 8576 10412 8628 10464
rect 9312 10412 9364 10464
rect 12072 10480 12124 10532
rect 1550 10310 1602 10362
rect 1614 10310 1666 10362
rect 1678 10310 1730 10362
rect 1742 10310 1794 10362
rect 1806 10310 1858 10362
rect 3550 10310 3602 10362
rect 3614 10310 3666 10362
rect 3678 10310 3730 10362
rect 3742 10310 3794 10362
rect 3806 10310 3858 10362
rect 5550 10310 5602 10362
rect 5614 10310 5666 10362
rect 5678 10310 5730 10362
rect 5742 10310 5794 10362
rect 5806 10310 5858 10362
rect 7550 10310 7602 10362
rect 7614 10310 7666 10362
rect 7678 10310 7730 10362
rect 7742 10310 7794 10362
rect 7806 10310 7858 10362
rect 9550 10310 9602 10362
rect 9614 10310 9666 10362
rect 9678 10310 9730 10362
rect 9742 10310 9794 10362
rect 9806 10310 9858 10362
rect 11550 10310 11602 10362
rect 11614 10310 11666 10362
rect 11678 10310 11730 10362
rect 11742 10310 11794 10362
rect 11806 10310 11858 10362
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 11980 10208 12032 10260
rect 1492 10115 1544 10124
rect 1492 10081 1501 10115
rect 1501 10081 1535 10115
rect 1535 10081 1544 10115
rect 1492 10072 1544 10081
rect 1952 10115 2004 10124
rect 1952 10081 1961 10115
rect 1961 10081 1995 10115
rect 1995 10081 2004 10115
rect 1952 10072 2004 10081
rect 2688 10072 2740 10124
rect 3884 10004 3936 10056
rect 3332 9936 3384 9988
rect 4620 10004 4672 10056
rect 6920 10072 6972 10124
rect 8852 10072 8904 10124
rect 5908 9936 5960 9988
rect 8484 10004 8536 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 9772 10004 9824 10056
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 8944 9979 8996 9988
rect 8944 9945 8953 9979
rect 8953 9945 8987 9979
rect 8987 9945 8996 9979
rect 8944 9936 8996 9945
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 7288 9868 7340 9920
rect 8116 9911 8168 9920
rect 8116 9877 8125 9911
rect 8125 9877 8159 9911
rect 8159 9877 8168 9911
rect 8116 9868 8168 9877
rect 8668 9868 8720 9920
rect 11244 9936 11296 9988
rect 11336 9979 11388 9988
rect 11336 9945 11345 9979
rect 11345 9945 11379 9979
rect 11379 9945 11388 9979
rect 11336 9936 11388 9945
rect 9956 9868 10008 9920
rect 10784 9911 10836 9920
rect 10784 9877 10793 9911
rect 10793 9877 10827 9911
rect 10827 9877 10836 9911
rect 10784 9868 10836 9877
rect 11428 9868 11480 9920
rect 2250 9766 2302 9818
rect 2314 9766 2366 9818
rect 2378 9766 2430 9818
rect 2442 9766 2494 9818
rect 2506 9766 2558 9818
rect 4250 9766 4302 9818
rect 4314 9766 4366 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 6250 9766 6302 9818
rect 6314 9766 6366 9818
rect 6378 9766 6430 9818
rect 6442 9766 6494 9818
rect 6506 9766 6558 9818
rect 8250 9766 8302 9818
rect 8314 9766 8366 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 10250 9766 10302 9818
rect 10314 9766 10366 9818
rect 10378 9766 10430 9818
rect 10442 9766 10494 9818
rect 10506 9766 10558 9818
rect 2688 9664 2740 9716
rect 1492 9596 1544 9648
rect 3424 9596 3476 9648
rect 5448 9596 5500 9648
rect 6644 9596 6696 9648
rect 8944 9664 8996 9716
rect 9772 9639 9824 9648
rect 9772 9605 9781 9639
rect 9781 9605 9815 9639
rect 9815 9605 9824 9639
rect 9772 9596 9824 9605
rect 10048 9596 10100 9648
rect 10876 9596 10928 9648
rect 6920 9528 6972 9580
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 9312 9528 9364 9580
rect 1400 9460 1452 9512
rect 7012 9460 7064 9512
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 10968 9528 11020 9580
rect 12164 9528 12216 9580
rect 11152 9460 11204 9512
rect 9404 9392 9456 9444
rect 2136 9324 2188 9376
rect 3976 9324 4028 9376
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 4620 9324 4672 9376
rect 6092 9324 6144 9376
rect 7932 9324 7984 9376
rect 1550 9222 1602 9274
rect 1614 9222 1666 9274
rect 1678 9222 1730 9274
rect 1742 9222 1794 9274
rect 1806 9222 1858 9274
rect 3550 9222 3602 9274
rect 3614 9222 3666 9274
rect 3678 9222 3730 9274
rect 3742 9222 3794 9274
rect 3806 9222 3858 9274
rect 5550 9222 5602 9274
rect 5614 9222 5666 9274
rect 5678 9222 5730 9274
rect 5742 9222 5794 9274
rect 5806 9222 5858 9274
rect 7550 9222 7602 9274
rect 7614 9222 7666 9274
rect 7678 9222 7730 9274
rect 7742 9222 7794 9274
rect 7806 9222 7858 9274
rect 9550 9222 9602 9274
rect 9614 9222 9666 9274
rect 9678 9222 9730 9274
rect 9742 9222 9794 9274
rect 9806 9222 9858 9274
rect 11550 9222 11602 9274
rect 11614 9222 11666 9274
rect 11678 9222 11730 9274
rect 11742 9222 11794 9274
rect 11806 9222 11858 9274
rect 2872 9120 2924 9172
rect 848 9052 900 9104
rect 2136 9052 2188 9104
rect 5908 9120 5960 9172
rect 6092 9163 6144 9172
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 8668 9120 8720 9172
rect 1400 8984 1452 9036
rect 4068 8984 4120 9036
rect 7288 9027 7340 9036
rect 7288 8993 7297 9027
rect 7297 8993 7331 9027
rect 7331 8993 7340 9027
rect 7288 8984 7340 8993
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 9956 8984 10008 9036
rect 2044 8916 2096 8968
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 3976 8916 4028 8968
rect 2872 8848 2924 8900
rect 3332 8891 3384 8900
rect 3332 8857 3341 8891
rect 3341 8857 3375 8891
rect 3375 8857 3384 8891
rect 3332 8848 3384 8857
rect 3424 8848 3476 8900
rect 4620 8848 4672 8900
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 5908 8916 5960 8968
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 6736 8916 6788 8968
rect 6184 8891 6236 8900
rect 6184 8857 6193 8891
rect 6193 8857 6227 8891
rect 6227 8857 6236 8891
rect 6184 8848 6236 8857
rect 3240 8780 3292 8832
rect 5448 8780 5500 8832
rect 6000 8780 6052 8832
rect 7932 8848 7984 8900
rect 8024 8780 8076 8832
rect 9036 8848 9088 8900
rect 9496 8848 9548 8900
rect 9128 8780 9180 8832
rect 10048 8916 10100 8968
rect 9956 8848 10008 8900
rect 10876 8848 10928 8900
rect 9864 8780 9916 8832
rect 10692 8780 10744 8832
rect 11152 8780 11204 8832
rect 2250 8678 2302 8730
rect 2314 8678 2366 8730
rect 2378 8678 2430 8730
rect 2442 8678 2494 8730
rect 2506 8678 2558 8730
rect 4250 8678 4302 8730
rect 4314 8678 4366 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 6250 8678 6302 8730
rect 6314 8678 6366 8730
rect 6378 8678 6430 8730
rect 6442 8678 6494 8730
rect 6506 8678 6558 8730
rect 8250 8678 8302 8730
rect 8314 8678 8366 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 10250 8678 10302 8730
rect 10314 8678 10366 8730
rect 10378 8678 10430 8730
rect 10442 8678 10494 8730
rect 10506 8678 10558 8730
rect 2136 8576 2188 8628
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 2596 8576 2648 8628
rect 5356 8576 5408 8628
rect 8668 8576 8720 8628
rect 9588 8576 9640 8628
rect 1952 8508 2004 8560
rect 2412 8440 2464 8492
rect 3332 8508 3384 8560
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 6736 8440 6788 8492
rect 8760 8508 8812 8560
rect 10048 8576 10100 8628
rect 10784 8576 10836 8628
rect 11244 8576 11296 8628
rect 9864 8508 9916 8560
rect 10140 8551 10192 8560
rect 10140 8517 10149 8551
rect 10149 8517 10183 8551
rect 10183 8517 10192 8551
rect 10140 8508 10192 8517
rect 2044 8415 2096 8424
rect 2044 8381 2053 8415
rect 2053 8381 2087 8415
rect 2087 8381 2096 8415
rect 2044 8372 2096 8381
rect 2320 8372 2372 8424
rect 2688 8372 2740 8424
rect 3424 8372 3476 8424
rect 848 8304 900 8356
rect 1952 8304 2004 8356
rect 7932 8440 7984 8492
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 9588 8440 9640 8492
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 10048 8372 10100 8424
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 11152 8508 11204 8560
rect 11428 8440 11480 8492
rect 12072 8576 12124 8628
rect 9588 8304 9640 8356
rect 12164 8372 12216 8424
rect 3332 8236 3384 8288
rect 6000 8236 6052 8288
rect 7288 8236 7340 8288
rect 12072 8304 12124 8356
rect 10324 8279 10376 8288
rect 10324 8245 10333 8279
rect 10333 8245 10367 8279
rect 10367 8245 10376 8279
rect 10324 8236 10376 8245
rect 1550 8134 1602 8186
rect 1614 8134 1666 8186
rect 1678 8134 1730 8186
rect 1742 8134 1794 8186
rect 1806 8134 1858 8186
rect 3550 8134 3602 8186
rect 3614 8134 3666 8186
rect 3678 8134 3730 8186
rect 3742 8134 3794 8186
rect 3806 8134 3858 8186
rect 5550 8134 5602 8186
rect 5614 8134 5666 8186
rect 5678 8134 5730 8186
rect 5742 8134 5794 8186
rect 5806 8134 5858 8186
rect 7550 8134 7602 8186
rect 7614 8134 7666 8186
rect 7678 8134 7730 8186
rect 7742 8134 7794 8186
rect 7806 8134 7858 8186
rect 9550 8134 9602 8186
rect 9614 8134 9666 8186
rect 9678 8134 9730 8186
rect 9742 8134 9794 8186
rect 9806 8134 9858 8186
rect 11550 8134 11602 8186
rect 11614 8134 11666 8186
rect 11678 8134 11730 8186
rect 11742 8134 11794 8186
rect 11806 8134 11858 8186
rect 6644 8075 6696 8084
rect 6644 8041 6653 8075
rect 6653 8041 6687 8075
rect 6687 8041 6696 8075
rect 6644 8032 6696 8041
rect 8852 8032 8904 8084
rect 9956 8032 10008 8084
rect 10876 8032 10928 8084
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 11888 8032 11940 8084
rect 2320 8007 2372 8016
rect 2320 7973 2329 8007
rect 2329 7973 2363 8007
rect 2363 7973 2372 8007
rect 2320 7964 2372 7973
rect 9036 7964 9088 8016
rect 9220 7964 9272 8016
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 2044 7828 2096 7880
rect 2136 7760 2188 7812
rect 2596 7803 2648 7812
rect 2596 7769 2605 7803
rect 2605 7769 2639 7803
rect 2639 7769 2648 7803
rect 2596 7760 2648 7769
rect 4160 7828 4212 7880
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 8760 7828 8812 7880
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 9956 7896 10008 7948
rect 10324 7896 10376 7948
rect 9496 7828 9548 7880
rect 10048 7828 10100 7880
rect 11152 7964 11204 8016
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 11336 7828 11388 7880
rect 848 7692 900 7744
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 3424 7692 3476 7744
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 2250 7590 2302 7642
rect 2314 7590 2366 7642
rect 2378 7590 2430 7642
rect 2442 7590 2494 7642
rect 2506 7590 2558 7642
rect 4250 7590 4302 7642
rect 4314 7590 4366 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 6250 7590 6302 7642
rect 6314 7590 6366 7642
rect 6378 7590 6430 7642
rect 6442 7590 6494 7642
rect 6506 7590 6558 7642
rect 8250 7590 8302 7642
rect 8314 7590 8366 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 10250 7590 10302 7642
rect 10314 7590 10366 7642
rect 10378 7590 10430 7642
rect 10442 7590 10494 7642
rect 10506 7590 10558 7642
rect 2688 7488 2740 7540
rect 8668 7488 8720 7540
rect 1400 7352 1452 7404
rect 3976 7352 4028 7404
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 8668 7352 8720 7404
rect 1860 7284 1912 7336
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 9036 7284 9088 7336
rect 10968 7352 11020 7404
rect 11980 7284 12032 7336
rect 8300 7216 8352 7268
rect 11244 7148 11296 7200
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 11888 7148 11940 7200
rect 1550 7046 1602 7098
rect 1614 7046 1666 7098
rect 1678 7046 1730 7098
rect 1742 7046 1794 7098
rect 1806 7046 1858 7098
rect 3550 7046 3602 7098
rect 3614 7046 3666 7098
rect 3678 7046 3730 7098
rect 3742 7046 3794 7098
rect 3806 7046 3858 7098
rect 5550 7046 5602 7098
rect 5614 7046 5666 7098
rect 5678 7046 5730 7098
rect 5742 7046 5794 7098
rect 5806 7046 5858 7098
rect 7550 7046 7602 7098
rect 7614 7046 7666 7098
rect 7678 7046 7730 7098
rect 7742 7046 7794 7098
rect 7806 7046 7858 7098
rect 9550 7046 9602 7098
rect 9614 7046 9666 7098
rect 9678 7046 9730 7098
rect 9742 7046 9794 7098
rect 9806 7046 9858 7098
rect 11550 7046 11602 7098
rect 11614 7046 11666 7098
rect 11678 7046 11730 7098
rect 11742 7046 11794 7098
rect 11806 7046 11858 7098
rect 1952 6944 2004 6996
rect 7288 6944 7340 6996
rect 2044 6808 2096 6860
rect 6920 6808 6972 6860
rect 7932 6808 7984 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9956 6876 10008 6928
rect 10784 6808 10836 6860
rect 8300 6740 8352 6792
rect 8852 6740 8904 6792
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 2044 6672 2096 6724
rect 10140 6672 10192 6724
rect 11244 6672 11296 6724
rect 11980 6604 12032 6656
rect 2250 6502 2302 6554
rect 2314 6502 2366 6554
rect 2378 6502 2430 6554
rect 2442 6502 2494 6554
rect 2506 6502 2558 6554
rect 4250 6502 4302 6554
rect 4314 6502 4366 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 6250 6502 6302 6554
rect 6314 6502 6366 6554
rect 6378 6502 6430 6554
rect 6442 6502 6494 6554
rect 6506 6502 6558 6554
rect 8250 6502 8302 6554
rect 8314 6502 8366 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 10250 6502 10302 6554
rect 10314 6502 10366 6554
rect 10378 6502 10430 6554
rect 10442 6502 10494 6554
rect 10506 6502 10558 6554
rect 8852 6443 8904 6452
rect 8852 6409 8861 6443
rect 8861 6409 8895 6443
rect 8895 6409 8904 6443
rect 8852 6400 8904 6409
rect 1952 6375 2004 6384
rect 1952 6341 1961 6375
rect 1961 6341 1995 6375
rect 1995 6341 2004 6375
rect 1952 6332 2004 6341
rect 2044 6332 2096 6384
rect 3332 6332 3384 6384
rect 4896 6375 4948 6384
rect 848 6060 900 6112
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 4896 6341 4905 6375
rect 4905 6341 4939 6375
rect 4939 6341 4948 6375
rect 4896 6332 4948 6341
rect 5080 6375 5132 6384
rect 5080 6341 5105 6375
rect 5105 6341 5132 6375
rect 5080 6332 5132 6341
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 9956 6332 10008 6384
rect 10600 6332 10652 6384
rect 11428 6264 11480 6316
rect 2596 6196 2648 6248
rect 2964 6128 3016 6180
rect 3056 6171 3108 6180
rect 3056 6137 3065 6171
rect 3065 6137 3099 6171
rect 3099 6137 3108 6171
rect 3056 6128 3108 6137
rect 9404 6239 9456 6248
rect 9404 6205 9413 6239
rect 9413 6205 9447 6239
rect 9447 6205 9456 6239
rect 9404 6196 9456 6205
rect 2596 6060 2648 6112
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 3424 6060 3476 6112
rect 4160 6060 4212 6112
rect 11152 6128 11204 6180
rect 5356 6060 5408 6112
rect 10048 6060 10100 6112
rect 11244 6060 11296 6112
rect 12164 6060 12216 6112
rect 1550 5958 1602 6010
rect 1614 5958 1666 6010
rect 1678 5958 1730 6010
rect 1742 5958 1794 6010
rect 1806 5958 1858 6010
rect 3550 5958 3602 6010
rect 3614 5958 3666 6010
rect 3678 5958 3730 6010
rect 3742 5958 3794 6010
rect 3806 5958 3858 6010
rect 5550 5958 5602 6010
rect 5614 5958 5666 6010
rect 5678 5958 5730 6010
rect 5742 5958 5794 6010
rect 5806 5958 5858 6010
rect 7550 5958 7602 6010
rect 7614 5958 7666 6010
rect 7678 5958 7730 6010
rect 7742 5958 7794 6010
rect 7806 5958 7858 6010
rect 9550 5958 9602 6010
rect 9614 5958 9666 6010
rect 9678 5958 9730 6010
rect 9742 5958 9794 6010
rect 9806 5958 9858 6010
rect 11550 5958 11602 6010
rect 11614 5958 11666 6010
rect 11678 5958 11730 6010
rect 11742 5958 11794 6010
rect 11806 5958 11858 6010
rect 1952 5856 2004 5908
rect 2872 5856 2924 5908
rect 10048 5856 10100 5908
rect 9772 5788 9824 5840
rect 2872 5720 2924 5772
rect 3148 5720 3200 5772
rect 848 5516 900 5568
rect 4160 5652 4212 5704
rect 2136 5627 2188 5636
rect 2136 5593 2145 5627
rect 2145 5593 2179 5627
rect 2179 5593 2188 5627
rect 2136 5584 2188 5593
rect 3424 5584 3476 5636
rect 7288 5652 7340 5704
rect 8576 5720 8628 5772
rect 9036 5720 9088 5772
rect 10692 5720 10744 5772
rect 10784 5720 10836 5772
rect 5908 5627 5960 5636
rect 5908 5593 5917 5627
rect 5917 5593 5951 5627
rect 5951 5593 5960 5627
rect 5908 5584 5960 5593
rect 1952 5516 2004 5568
rect 2964 5516 3016 5568
rect 3884 5516 3936 5568
rect 5448 5516 5500 5568
rect 7288 5516 7340 5568
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 8116 5584 8168 5636
rect 9956 5584 10008 5636
rect 11244 5720 11296 5772
rect 10968 5584 11020 5636
rect 11336 5584 11388 5636
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 11796 5559 11848 5568
rect 11796 5525 11805 5559
rect 11805 5525 11839 5559
rect 11839 5525 11848 5559
rect 11796 5516 11848 5525
rect 2250 5414 2302 5466
rect 2314 5414 2366 5466
rect 2378 5414 2430 5466
rect 2442 5414 2494 5466
rect 2506 5414 2558 5466
rect 4250 5414 4302 5466
rect 4314 5414 4366 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 6250 5414 6302 5466
rect 6314 5414 6366 5466
rect 6378 5414 6430 5466
rect 6442 5414 6494 5466
rect 6506 5414 6558 5466
rect 8250 5414 8302 5466
rect 8314 5414 8366 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 10250 5414 10302 5466
rect 10314 5414 10366 5466
rect 10378 5414 10430 5466
rect 10442 5414 10494 5466
rect 10506 5414 10558 5466
rect 3884 5355 3936 5364
rect 3884 5321 3893 5355
rect 3893 5321 3927 5355
rect 3927 5321 3936 5355
rect 3884 5312 3936 5321
rect 4068 5312 4120 5364
rect 5080 5312 5132 5364
rect 5908 5312 5960 5364
rect 9496 5312 9548 5364
rect 3332 5244 3384 5296
rect 2872 5176 2924 5228
rect 3424 5176 3476 5228
rect 4620 5176 4672 5228
rect 4896 5176 4948 5228
rect 5908 5176 5960 5228
rect 6920 5244 6972 5296
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 7472 5244 7524 5296
rect 7104 5176 7156 5228
rect 8116 5244 8168 5296
rect 8668 5244 8720 5296
rect 10140 5312 10192 5364
rect 10600 5312 10652 5364
rect 10784 5287 10836 5296
rect 10784 5253 10811 5287
rect 10811 5253 10836 5287
rect 10784 5244 10836 5253
rect 11244 5312 11296 5364
rect 11152 5244 11204 5296
rect 11796 5244 11848 5296
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 1860 5108 1912 5160
rect 2136 5108 2188 5160
rect 8944 5108 8996 5160
rect 10140 5176 10192 5228
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 11060 5176 11112 5228
rect 12164 5176 12216 5228
rect 10692 5040 10744 5092
rect 10048 4972 10100 5024
rect 11060 4972 11112 5024
rect 11336 4972 11388 5024
rect 11980 5040 12032 5092
rect 1550 4870 1602 4922
rect 1614 4870 1666 4922
rect 1678 4870 1730 4922
rect 1742 4870 1794 4922
rect 1806 4870 1858 4922
rect 3550 4870 3602 4922
rect 3614 4870 3666 4922
rect 3678 4870 3730 4922
rect 3742 4870 3794 4922
rect 3806 4870 3858 4922
rect 5550 4870 5602 4922
rect 5614 4870 5666 4922
rect 5678 4870 5730 4922
rect 5742 4870 5794 4922
rect 5806 4870 5858 4922
rect 7550 4870 7602 4922
rect 7614 4870 7666 4922
rect 7678 4870 7730 4922
rect 7742 4870 7794 4922
rect 7806 4870 7858 4922
rect 9550 4870 9602 4922
rect 9614 4870 9666 4922
rect 9678 4870 9730 4922
rect 9742 4870 9794 4922
rect 9806 4870 9858 4922
rect 11550 4870 11602 4922
rect 11614 4870 11666 4922
rect 11678 4870 11730 4922
rect 11742 4870 11794 4922
rect 11806 4870 11858 4922
rect 3056 4811 3108 4820
rect 3056 4777 3065 4811
rect 3065 4777 3099 4811
rect 3099 4777 3108 4811
rect 3056 4768 3108 4777
rect 3332 4700 3384 4752
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 3884 4632 3936 4684
rect 6000 4632 6052 4684
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 2596 4496 2648 4548
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 7380 4768 7432 4820
rect 9956 4768 10008 4820
rect 10784 4768 10836 4820
rect 11888 4768 11940 4820
rect 9496 4700 9548 4752
rect 12072 4700 12124 4752
rect 7104 4632 7156 4684
rect 8024 4632 8076 4684
rect 11152 4632 11204 4684
rect 3240 4428 3292 4480
rect 4160 4428 4212 4480
rect 6644 4496 6696 4548
rect 8116 4564 8168 4616
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 9404 4496 9456 4548
rect 10232 4428 10284 4480
rect 10692 4428 10744 4480
rect 11152 4539 11204 4548
rect 11152 4505 11161 4539
rect 11161 4505 11195 4539
rect 11195 4505 11204 4539
rect 11152 4496 11204 4505
rect 11336 4428 11388 4480
rect 2250 4326 2302 4378
rect 2314 4326 2366 4378
rect 2378 4326 2430 4378
rect 2442 4326 2494 4378
rect 2506 4326 2558 4378
rect 4250 4326 4302 4378
rect 4314 4326 4366 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 6250 4326 6302 4378
rect 6314 4326 6366 4378
rect 6378 4326 6430 4378
rect 6442 4326 6494 4378
rect 6506 4326 6558 4378
rect 8250 4326 8302 4378
rect 8314 4326 8366 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 10250 4326 10302 4378
rect 10314 4326 10366 4378
rect 10378 4326 10430 4378
rect 10442 4326 10494 4378
rect 10506 4326 10558 4378
rect 5724 4224 5776 4276
rect 7288 4224 7340 4276
rect 9404 4267 9456 4276
rect 6092 4156 6144 4208
rect 4160 4088 4212 4140
rect 6920 4156 6972 4208
rect 3240 4020 3292 4072
rect 3424 4063 3476 4072
rect 3424 4029 3433 4063
rect 3433 4029 3467 4063
rect 3467 4029 3476 4063
rect 3424 4020 3476 4029
rect 3976 4020 4028 4072
rect 4620 4020 4672 4072
rect 3884 3952 3936 4004
rect 4252 3952 4304 4004
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 8024 4131 8076 4140
rect 8024 4097 8033 4131
rect 8033 4097 8067 4131
rect 8067 4097 8076 4131
rect 8024 4088 8076 4097
rect 9404 4233 9413 4267
rect 9413 4233 9447 4267
rect 9447 4233 9456 4267
rect 9404 4224 9456 4233
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 10416 4224 10468 4276
rect 6184 3995 6236 4004
rect 6184 3961 6193 3995
rect 6193 3961 6227 3995
rect 6227 3961 6236 3995
rect 8484 4020 8536 4072
rect 9496 4088 9548 4140
rect 11152 4131 11204 4140
rect 11152 4097 11161 4131
rect 11161 4097 11195 4131
rect 11195 4097 11204 4131
rect 11152 4088 11204 4097
rect 10140 4020 10192 4072
rect 10416 4063 10468 4072
rect 10416 4029 10425 4063
rect 10425 4029 10459 4063
rect 10459 4029 10468 4063
rect 10416 4020 10468 4029
rect 12164 4020 12216 4072
rect 6184 3952 6236 3961
rect 11796 3995 11848 4004
rect 11796 3961 11805 3995
rect 11805 3961 11839 3995
rect 11839 3961 11848 3995
rect 11796 3952 11848 3961
rect 2688 3927 2740 3936
rect 2688 3893 2697 3927
rect 2697 3893 2731 3927
rect 2731 3893 2740 3927
rect 2688 3884 2740 3893
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 5172 3884 5224 3936
rect 5908 3884 5960 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 9404 3884 9456 3936
rect 1550 3782 1602 3834
rect 1614 3782 1666 3834
rect 1678 3782 1730 3834
rect 1742 3782 1794 3834
rect 1806 3782 1858 3834
rect 3550 3782 3602 3834
rect 3614 3782 3666 3834
rect 3678 3782 3730 3834
rect 3742 3782 3794 3834
rect 3806 3782 3858 3834
rect 5550 3782 5602 3834
rect 5614 3782 5666 3834
rect 5678 3782 5730 3834
rect 5742 3782 5794 3834
rect 5806 3782 5858 3834
rect 7550 3782 7602 3834
rect 7614 3782 7666 3834
rect 7678 3782 7730 3834
rect 7742 3782 7794 3834
rect 7806 3782 7858 3834
rect 9550 3782 9602 3834
rect 9614 3782 9666 3834
rect 9678 3782 9730 3834
rect 9742 3782 9794 3834
rect 9806 3782 9858 3834
rect 11550 3782 11602 3834
rect 11614 3782 11666 3834
rect 11678 3782 11730 3834
rect 11742 3782 11794 3834
rect 11806 3782 11858 3834
rect 1952 3680 2004 3732
rect 6000 3680 6052 3732
rect 8116 3680 8168 3732
rect 4160 3587 4212 3596
rect 4160 3553 4169 3587
rect 4169 3553 4203 3587
rect 4203 3553 4212 3587
rect 4160 3544 4212 3553
rect 5448 3544 5500 3596
rect 6276 3544 6328 3596
rect 6736 3544 6788 3596
rect 10692 3680 10744 3732
rect 11152 3680 11204 3732
rect 2136 3451 2188 3460
rect 2136 3417 2145 3451
rect 2145 3417 2179 3451
rect 2179 3417 2188 3451
rect 2136 3408 2188 3417
rect 7380 3476 7432 3528
rect 8024 3476 8076 3528
rect 8484 3476 8536 3528
rect 9404 3476 9456 3528
rect 4160 3408 4212 3460
rect 4712 3408 4764 3460
rect 5172 3408 5224 3460
rect 3424 3340 3476 3392
rect 5816 3340 5868 3392
rect 6184 3408 6236 3460
rect 6092 3340 6144 3392
rect 6368 3340 6420 3392
rect 9956 3544 10008 3596
rect 10416 3544 10468 3596
rect 10968 3544 11020 3596
rect 9864 3408 9916 3460
rect 10048 3408 10100 3460
rect 10692 3408 10744 3460
rect 7656 3340 7708 3392
rect 11796 3383 11848 3392
rect 11796 3349 11805 3383
rect 11805 3349 11839 3383
rect 11839 3349 11848 3383
rect 11796 3340 11848 3349
rect 2250 3238 2302 3290
rect 2314 3238 2366 3290
rect 2378 3238 2430 3290
rect 2442 3238 2494 3290
rect 2506 3238 2558 3290
rect 4250 3238 4302 3290
rect 4314 3238 4366 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 6250 3238 6302 3290
rect 6314 3238 6366 3290
rect 6378 3238 6430 3290
rect 6442 3238 6494 3290
rect 6506 3238 6558 3290
rect 8250 3238 8302 3290
rect 8314 3238 8366 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 10250 3238 10302 3290
rect 10314 3238 10366 3290
rect 10378 3238 10430 3290
rect 10442 3238 10494 3290
rect 10506 3238 10558 3290
rect 2688 3136 2740 3188
rect 1952 3068 2004 3120
rect 4620 3179 4672 3188
rect 4620 3145 4629 3179
rect 4629 3145 4663 3179
rect 4663 3145 4672 3179
rect 4620 3136 4672 3145
rect 5356 3136 5408 3188
rect 2780 3000 2832 3052
rect 4436 3068 4488 3120
rect 5908 3068 5960 3120
rect 6000 3068 6052 3120
rect 6828 3136 6880 3188
rect 7104 3068 7156 3120
rect 7564 3068 7616 3120
rect 2136 2932 2188 2984
rect 2596 2932 2648 2984
rect 4712 2932 4764 2984
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 6736 3000 6788 3052
rect 11428 3136 11480 3188
rect 9036 3000 9088 3052
rect 9956 3068 10008 3120
rect 11244 3068 11296 3120
rect 11980 3000 12032 3052
rect 7932 2975 7984 2984
rect 7932 2941 7941 2975
rect 7941 2941 7975 2975
rect 7975 2941 7984 2975
rect 7932 2932 7984 2941
rect 9864 2975 9916 2984
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 7012 2864 7064 2916
rect 10968 2864 11020 2916
rect 6092 2796 6144 2848
rect 6368 2796 6420 2848
rect 6920 2796 6972 2848
rect 9956 2796 10008 2848
rect 1550 2694 1602 2746
rect 1614 2694 1666 2746
rect 1678 2694 1730 2746
rect 1742 2694 1794 2746
rect 1806 2694 1858 2746
rect 3550 2694 3602 2746
rect 3614 2694 3666 2746
rect 3678 2694 3730 2746
rect 3742 2694 3794 2746
rect 3806 2694 3858 2746
rect 5550 2694 5602 2746
rect 5614 2694 5666 2746
rect 5678 2694 5730 2746
rect 5742 2694 5794 2746
rect 5806 2694 5858 2746
rect 7550 2694 7602 2746
rect 7614 2694 7666 2746
rect 7678 2694 7730 2746
rect 7742 2694 7794 2746
rect 7806 2694 7858 2746
rect 9550 2694 9602 2746
rect 9614 2694 9666 2746
rect 9678 2694 9730 2746
rect 9742 2694 9794 2746
rect 9806 2694 9858 2746
rect 11550 2694 11602 2746
rect 11614 2694 11666 2746
rect 11678 2694 11730 2746
rect 11742 2694 11794 2746
rect 11806 2694 11858 2746
rect 4436 2635 4488 2644
rect 4436 2601 4445 2635
rect 4445 2601 4479 2635
rect 4479 2601 4488 2635
rect 4436 2592 4488 2601
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 7380 2592 7432 2644
rect 7932 2592 7984 2644
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 10692 2592 10744 2644
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 11980 2592 12032 2644
rect 6920 2524 6972 2576
rect 3424 2388 3476 2440
rect 4620 2456 4672 2508
rect 6000 2456 6052 2508
rect 4160 2320 4212 2372
rect 6736 2388 6788 2440
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 7288 2388 7340 2440
rect 8024 2388 8076 2440
rect 9220 2456 9272 2508
rect 9956 2499 10008 2508
rect 9956 2465 9965 2499
rect 9965 2465 9999 2499
rect 9999 2465 10008 2499
rect 9956 2456 10008 2465
rect 11060 2431 11112 2440
rect 11060 2397 11069 2431
rect 11069 2397 11103 2431
rect 11103 2397 11112 2431
rect 11060 2388 11112 2397
rect 3240 2252 3292 2304
rect 3884 2252 3936 2304
rect 5816 2252 5868 2304
rect 6644 2295 6696 2304
rect 6644 2261 6653 2295
rect 6653 2261 6687 2295
rect 6687 2261 6696 2295
rect 6644 2252 6696 2261
rect 7104 2252 7156 2304
rect 7748 2252 7800 2304
rect 9036 2252 9088 2304
rect 2250 2150 2302 2202
rect 2314 2150 2366 2202
rect 2378 2150 2430 2202
rect 2442 2150 2494 2202
rect 2506 2150 2558 2202
rect 4250 2150 4302 2202
rect 4314 2150 4366 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 6250 2150 6302 2202
rect 6314 2150 6366 2202
rect 6378 2150 6430 2202
rect 6442 2150 6494 2202
rect 6506 2150 6558 2202
rect 8250 2150 8302 2202
rect 8314 2150 8366 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 10250 2150 10302 2202
rect 10314 2150 10366 2202
rect 10378 2150 10430 2202
rect 10442 2150 10494 2202
rect 10506 2150 10558 2202
<< metal2 >>
rect 4526 14906 4582 15551
rect 5170 14906 5226 15551
rect 4526 14878 4660 14906
rect 4526 14751 4582 14878
rect 2250 13084 2558 13093
rect 2250 13082 2256 13084
rect 2312 13082 2336 13084
rect 2392 13082 2416 13084
rect 2472 13082 2496 13084
rect 2552 13082 2558 13084
rect 2312 13030 2314 13082
rect 2494 13030 2496 13082
rect 2250 13028 2256 13030
rect 2312 13028 2336 13030
rect 2392 13028 2416 13030
rect 2472 13028 2496 13030
rect 2552 13028 2558 13030
rect 2250 13019 2558 13028
rect 4250 13084 4558 13093
rect 4250 13082 4256 13084
rect 4312 13082 4336 13084
rect 4392 13082 4416 13084
rect 4472 13082 4496 13084
rect 4552 13082 4558 13084
rect 4312 13030 4314 13082
rect 4494 13030 4496 13082
rect 4250 13028 4256 13030
rect 4312 13028 4336 13030
rect 4392 13028 4416 13030
rect 4472 13028 4496 13030
rect 4552 13028 4558 13030
rect 4250 13019 4558 13028
rect 4632 12986 4660 14878
rect 5000 14878 5226 14906
rect 5000 12986 5028 14878
rect 5170 14751 5226 14878
rect 5814 14906 5870 15551
rect 6458 14906 6514 15551
rect 5814 14878 6132 14906
rect 5814 14751 5870 14878
rect 6104 12986 6132 14878
rect 6458 14878 6776 14906
rect 6458 14751 6514 14878
rect 6250 13084 6558 13093
rect 6250 13082 6256 13084
rect 6312 13082 6336 13084
rect 6392 13082 6416 13084
rect 6472 13082 6496 13084
rect 6552 13082 6558 13084
rect 6312 13030 6314 13082
rect 6494 13030 6496 13082
rect 6250 13028 6256 13030
rect 6312 13028 6336 13030
rect 6392 13028 6416 13030
rect 6472 13028 6496 13030
rect 6552 13028 6558 13030
rect 6250 13019 6558 13028
rect 6748 12986 6776 14878
rect 8250 13084 8558 13093
rect 8250 13082 8256 13084
rect 8312 13082 8336 13084
rect 8392 13082 8416 13084
rect 8472 13082 8496 13084
rect 8552 13082 8558 13084
rect 8312 13030 8314 13082
rect 8494 13030 8496 13082
rect 8250 13028 8256 13030
rect 8312 13028 8336 13030
rect 8392 13028 8416 13030
rect 8472 13028 8496 13030
rect 8552 13028 8558 13030
rect 8250 13019 8558 13028
rect 10250 13084 10558 13093
rect 10250 13082 10256 13084
rect 10312 13082 10336 13084
rect 10392 13082 10416 13084
rect 10472 13082 10496 13084
rect 10552 13082 10558 13084
rect 10312 13030 10314 13082
rect 10494 13030 10496 13082
rect 10250 13028 10256 13030
rect 10312 13028 10336 13030
rect 10392 13028 10416 13030
rect 10472 13028 10496 13030
rect 10552 13028 10558 13030
rect 10250 13019 10558 13028
rect 10782 13016 10838 13025
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6736 12980 6788 12986
rect 10782 12951 10838 12960
rect 6736 12922 6788 12928
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 1550 12540 1858 12549
rect 1550 12538 1556 12540
rect 1612 12538 1636 12540
rect 1692 12538 1716 12540
rect 1772 12538 1796 12540
rect 1852 12538 1858 12540
rect 1612 12486 1614 12538
rect 1794 12486 1796 12538
rect 1550 12484 1556 12486
rect 1612 12484 1636 12486
rect 1692 12484 1716 12486
rect 1772 12484 1796 12486
rect 1852 12484 1858 12486
rect 1550 12475 1858 12484
rect 3550 12540 3858 12549
rect 3550 12538 3556 12540
rect 3612 12538 3636 12540
rect 3692 12538 3716 12540
rect 3772 12538 3796 12540
rect 3852 12538 3858 12540
rect 3612 12486 3614 12538
rect 3794 12486 3796 12538
rect 3550 12484 3556 12486
rect 3612 12484 3636 12486
rect 3692 12484 3716 12486
rect 3772 12484 3796 12486
rect 3852 12484 3858 12486
rect 3550 12475 3858 12484
rect 5184 12306 5212 12718
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 2250 11996 2558 12005
rect 2250 11994 2256 11996
rect 2312 11994 2336 11996
rect 2392 11994 2416 11996
rect 2472 11994 2496 11996
rect 2552 11994 2558 11996
rect 2312 11942 2314 11994
rect 2494 11942 2496 11994
rect 2250 11940 2256 11942
rect 2312 11940 2336 11942
rect 2392 11940 2416 11942
rect 2472 11940 2496 11942
rect 2552 11940 2558 11942
rect 2250 11931 2558 11940
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 1550 11452 1858 11461
rect 1550 11450 1556 11452
rect 1612 11450 1636 11452
rect 1692 11450 1716 11452
rect 1772 11450 1796 11452
rect 1852 11450 1858 11452
rect 1612 11398 1614 11450
rect 1794 11398 1796 11450
rect 1550 11396 1556 11398
rect 1612 11396 1636 11398
rect 1692 11396 1716 11398
rect 1772 11396 1796 11398
rect 1852 11396 1858 11398
rect 1550 11387 1858 11396
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 848 10464 900 10470
rect 848 10406 900 10412
rect 860 9489 888 10406
rect 1550 10364 1858 10373
rect 1550 10362 1556 10364
rect 1612 10362 1636 10364
rect 1692 10362 1716 10364
rect 1772 10362 1796 10364
rect 1852 10362 1858 10364
rect 1612 10310 1614 10362
rect 1794 10310 1796 10362
rect 1550 10308 1556 10310
rect 1612 10308 1636 10310
rect 1692 10308 1716 10310
rect 1772 10308 1796 10310
rect 1852 10308 1858 10310
rect 1550 10299 1858 10308
rect 1964 10130 1992 10950
rect 2250 10908 2558 10917
rect 2250 10906 2256 10908
rect 2312 10906 2336 10908
rect 2392 10906 2416 10908
rect 2472 10906 2496 10908
rect 2552 10906 2558 10908
rect 2312 10854 2314 10906
rect 2494 10854 2496 10906
rect 2250 10852 2256 10854
rect 2312 10852 2336 10854
rect 2392 10852 2416 10854
rect 2472 10852 2496 10854
rect 2552 10852 2558 10854
rect 2250 10843 2558 10852
rect 3068 10742 3096 11630
rect 3550 11452 3858 11461
rect 3550 11450 3556 11452
rect 3612 11450 3636 11452
rect 3692 11450 3716 11452
rect 3772 11450 3796 11452
rect 3852 11450 3858 11452
rect 3612 11398 3614 11450
rect 3794 11398 3796 11450
rect 3550 11396 3556 11398
rect 3612 11396 3636 11398
rect 3692 11396 3716 11398
rect 3772 11396 3796 11398
rect 3852 11396 3858 11398
rect 3550 11387 3858 11396
rect 3056 10736 3108 10742
rect 3056 10678 3108 10684
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2700 10130 2728 10610
rect 3550 10364 3858 10373
rect 3550 10362 3556 10364
rect 3612 10362 3636 10364
rect 3692 10362 3716 10364
rect 3772 10362 3796 10364
rect 3852 10362 3858 10364
rect 3612 10310 3614 10362
rect 3794 10310 3796 10362
rect 3550 10308 3556 10310
rect 3612 10308 3636 10310
rect 3692 10308 3716 10310
rect 3772 10308 3796 10310
rect 3852 10308 3858 10310
rect 3550 10299 3858 10308
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 1504 9654 1532 10066
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1400 9512 1452 9518
rect 846 9480 902 9489
rect 1400 9454 1452 9460
rect 846 9415 902 9424
rect 848 9104 900 9110
rect 846 9072 848 9081
rect 900 9072 902 9081
rect 1412 9042 1440 9454
rect 1550 9276 1858 9285
rect 1550 9274 1556 9276
rect 1612 9274 1636 9276
rect 1692 9274 1716 9276
rect 1772 9274 1796 9276
rect 1852 9274 1858 9276
rect 1612 9222 1614 9274
rect 1794 9222 1796 9274
rect 1550 9220 1556 9222
rect 1612 9220 1636 9222
rect 1692 9220 1716 9222
rect 1772 9220 1796 9222
rect 1852 9220 1858 9222
rect 1550 9211 1858 9220
rect 846 9007 902 9016
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 848 8356 900 8362
rect 848 8298 900 8304
rect 860 8129 888 8298
rect 846 8120 902 8129
rect 846 8055 902 8064
rect 848 7744 900 7750
rect 846 7712 848 7721
rect 900 7712 902 7721
rect 846 7647 902 7656
rect 1412 7410 1440 8978
rect 1964 8566 1992 10066
rect 2250 9820 2558 9829
rect 2250 9818 2256 9820
rect 2312 9818 2336 9820
rect 2392 9818 2416 9820
rect 2472 9818 2496 9820
rect 2552 9818 2558 9820
rect 2312 9766 2314 9818
rect 2494 9766 2496 9818
rect 2250 9764 2256 9766
rect 2312 9764 2336 9766
rect 2392 9764 2416 9766
rect 2472 9764 2496 9766
rect 2552 9764 2558 9766
rect 2250 9755 2558 9764
rect 2700 9722 2728 10066
rect 3896 10062 3924 12174
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4080 11830 4108 12038
rect 4172 11898 4200 12038
rect 4250 11996 4558 12005
rect 4250 11994 4256 11996
rect 4312 11994 4336 11996
rect 4392 11994 4416 11996
rect 4472 11994 4496 11996
rect 4552 11994 4558 11996
rect 4312 11942 4314 11994
rect 4494 11942 4496 11994
rect 4250 11940 4256 11942
rect 4312 11940 4336 11942
rect 4392 11940 4416 11942
rect 4472 11940 4496 11942
rect 4552 11940 4558 11942
rect 4250 11931 4558 11940
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 4158 11656 4214 11665
rect 5184 11626 5212 12242
rect 5276 12238 5304 12786
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5828 12730 5856 12786
rect 5460 12442 5488 12718
rect 5828 12702 5948 12730
rect 5550 12540 5858 12549
rect 5550 12538 5556 12540
rect 5612 12538 5636 12540
rect 5692 12538 5716 12540
rect 5772 12538 5796 12540
rect 5852 12538 5858 12540
rect 5612 12486 5614 12538
rect 5794 12486 5796 12538
rect 5550 12484 5556 12486
rect 5612 12484 5636 12486
rect 5692 12484 5716 12486
rect 5772 12484 5796 12486
rect 5852 12484 5858 12486
rect 5550 12475 5858 12484
rect 5920 12442 5948 12702
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 4158 11591 4214 11600
rect 5172 11620 5224 11626
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 11218 4016 11494
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3988 11014 4016 11154
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2148 9110 2176 9318
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2044 8968 2096 8974
rect 2148 8922 2176 9046
rect 2096 8916 2176 8922
rect 2044 8910 2176 8916
rect 2056 8894 2176 8910
rect 2148 8634 2176 8894
rect 2250 8732 2558 8741
rect 2250 8730 2256 8732
rect 2312 8730 2336 8732
rect 2392 8730 2416 8732
rect 2472 8730 2496 8732
rect 2552 8730 2558 8732
rect 2312 8678 2314 8730
rect 2494 8678 2496 8730
rect 2250 8676 2256 8678
rect 2312 8676 2336 8678
rect 2392 8676 2416 8678
rect 2472 8676 2496 8678
rect 2552 8676 2558 8678
rect 2250 8667 2558 8676
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1550 8188 1858 8197
rect 1550 8186 1556 8188
rect 1612 8186 1636 8188
rect 1692 8186 1716 8188
rect 1772 8186 1796 8188
rect 1852 8186 1858 8188
rect 1612 8134 1614 8186
rect 1794 8134 1796 8186
rect 1550 8132 1556 8134
rect 1612 8132 1636 8134
rect 1692 8132 1716 8134
rect 1772 8132 1796 8134
rect 1852 8132 1858 8134
rect 1550 8123 1858 8132
rect 1964 7562 1992 8298
rect 2056 7886 2084 8366
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2148 7818 2176 8570
rect 2424 8498 2452 8570
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2332 8022 2360 8366
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2608 7818 2636 8570
rect 2700 8430 2728 9658
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2884 8906 2912 9114
rect 3344 8906 3372 9930
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 9654 3464 9862
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 4080 9382 4108 10678
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3550 9276 3858 9285
rect 3550 9274 3556 9276
rect 3612 9274 3636 9276
rect 3692 9274 3716 9276
rect 3772 9274 3796 9276
rect 3852 9274 3858 9276
rect 3612 9222 3614 9274
rect 3794 9222 3796 9274
rect 3550 9220 3556 9222
rect 3612 9220 3636 9222
rect 3692 9220 3716 9222
rect 3772 9220 3796 9222
rect 3852 9220 3858 9222
rect 3550 9211 3858 9220
rect 3988 8974 4016 9318
rect 4080 9042 4108 9318
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 8498 3280 8774
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 3344 8294 3372 8502
rect 3436 8430 3464 8842
rect 3804 8498 3832 8910
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2250 7644 2558 7653
rect 2250 7642 2256 7644
rect 2312 7642 2336 7644
rect 2392 7642 2416 7644
rect 2472 7642 2496 7644
rect 2552 7642 2558 7644
rect 2312 7590 2314 7642
rect 2494 7590 2496 7642
rect 2250 7588 2256 7590
rect 2312 7588 2336 7590
rect 2392 7588 2416 7590
rect 2472 7588 2496 7590
rect 2552 7588 2558 7590
rect 2250 7579 2558 7588
rect 1964 7534 2084 7562
rect 2700 7546 2728 7686
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1860 7336 1912 7342
rect 1912 7296 1992 7324
rect 1860 7278 1912 7284
rect 1550 7100 1858 7109
rect 1550 7098 1556 7100
rect 1612 7098 1636 7100
rect 1692 7098 1716 7100
rect 1772 7098 1796 7100
rect 1852 7098 1858 7100
rect 1612 7046 1614 7098
rect 1794 7046 1796 7098
rect 1550 7044 1556 7046
rect 1612 7044 1636 7046
rect 1692 7044 1716 7046
rect 1772 7044 1796 7046
rect 1852 7044 1858 7046
rect 1550 7035 1858 7044
rect 1964 7002 1992 7296
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2056 6866 2084 7534
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 2056 6390 2084 6666
rect 2250 6556 2558 6565
rect 2250 6554 2256 6556
rect 2312 6554 2336 6556
rect 2392 6554 2416 6556
rect 2472 6554 2496 6556
rect 2552 6554 2558 6556
rect 2312 6502 2314 6554
rect 2494 6502 2496 6554
rect 2250 6500 2256 6502
rect 2312 6500 2336 6502
rect 2392 6500 2416 6502
rect 2472 6500 2496 6502
rect 2552 6500 2558 6502
rect 2250 6491 2558 6500
rect 3344 6390 3372 8230
rect 3550 8188 3858 8197
rect 3550 8186 3556 8188
rect 3612 8186 3636 8188
rect 3692 8186 3716 8188
rect 3772 8186 3796 8188
rect 3852 8186 3858 8188
rect 3612 8134 3614 8186
rect 3794 8134 3796 8186
rect 3550 8132 3556 8134
rect 3612 8132 3636 8134
rect 3692 8132 3716 8134
rect 3772 8132 3796 8134
rect 3852 8132 3858 8134
rect 3550 8123 3858 8132
rect 4172 7886 4200 11591
rect 5172 11562 5224 11568
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4250 10908 4558 10917
rect 4250 10906 4256 10908
rect 4312 10906 4336 10908
rect 4392 10906 4416 10908
rect 4472 10906 4496 10908
rect 4552 10906 4558 10908
rect 4312 10854 4314 10906
rect 4494 10854 4496 10906
rect 4250 10852 4256 10854
rect 4312 10852 4336 10854
rect 4392 10852 4416 10854
rect 4472 10852 4496 10854
rect 4552 10852 4558 10854
rect 4250 10843 4558 10852
rect 4632 10606 4660 11154
rect 5184 11150 5212 11562
rect 5276 11354 5304 12174
rect 5460 11898 5488 12378
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5920 11762 5948 12038
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5368 11558 5396 11698
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5276 11082 5304 11290
rect 5368 11286 5396 11494
rect 5460 11354 5488 11698
rect 6012 11694 6040 12786
rect 6656 12306 6684 12786
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6250 11996 6558 12005
rect 6250 11994 6256 11996
rect 6312 11994 6336 11996
rect 6392 11994 6416 11996
rect 6472 11994 6496 11996
rect 6552 11994 6558 11996
rect 6312 11942 6314 11994
rect 6494 11942 6496 11994
rect 6250 11940 6256 11942
rect 6312 11940 6336 11942
rect 6392 11940 6416 11942
rect 6472 11940 6496 11942
rect 6552 11940 6558 11942
rect 6250 11931 6558 11940
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5550 11452 5858 11461
rect 5550 11450 5556 11452
rect 5612 11450 5636 11452
rect 5692 11450 5716 11452
rect 5772 11450 5796 11452
rect 5852 11450 5858 11452
rect 5612 11398 5614 11450
rect 5794 11398 5796 11450
rect 5550 11396 5556 11398
rect 5612 11396 5636 11398
rect 5692 11396 5716 11398
rect 5772 11396 5796 11398
rect 5852 11396 5858 11398
rect 5550 11387 5858 11396
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 6012 11218 6040 11630
rect 6656 11626 6684 12242
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6104 11218 6132 11494
rect 6932 11354 6960 12174
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11830 7236 12038
rect 7196 11824 7248 11830
rect 7196 11766 7248 11772
rect 7392 11694 7420 12650
rect 7550 12540 7858 12549
rect 7550 12538 7556 12540
rect 7612 12538 7636 12540
rect 7692 12538 7716 12540
rect 7772 12538 7796 12540
rect 7852 12538 7858 12540
rect 7612 12486 7614 12538
rect 7794 12486 7796 12538
rect 7550 12484 7556 12486
rect 7612 12484 7636 12486
rect 7692 12484 7716 12486
rect 7772 12484 7796 12486
rect 7852 12484 7858 12486
rect 7550 12475 7858 12484
rect 9550 12540 9858 12549
rect 9550 12538 9556 12540
rect 9612 12538 9636 12540
rect 9692 12538 9716 12540
rect 9772 12538 9796 12540
rect 9852 12538 9858 12540
rect 9612 12486 9614 12538
rect 9794 12486 9796 12538
rect 9550 12484 9556 12486
rect 9612 12484 9636 12486
rect 9692 12484 9716 12486
rect 9772 12484 9796 12486
rect 9852 12484 9858 12486
rect 9550 12475 9858 12484
rect 9968 12238 9996 12786
rect 10060 12306 10088 12786
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 8250 11996 8558 12005
rect 8250 11994 8256 11996
rect 8312 11994 8336 11996
rect 8392 11994 8416 11996
rect 8472 11994 8496 11996
rect 8552 11994 8558 11996
rect 8312 11942 8314 11994
rect 8494 11942 8496 11994
rect 8250 11940 8256 11942
rect 8312 11940 8336 11942
rect 8392 11940 8416 11942
rect 8472 11940 8496 11942
rect 8552 11940 8558 11942
rect 8250 11931 8558 11940
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 7104 11552 7156 11558
rect 7024 11500 7104 11506
rect 7024 11494 7156 11500
rect 7024 11478 7144 11494
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 6012 10810 6040 11154
rect 6250 10908 6558 10917
rect 6250 10906 6256 10908
rect 6312 10906 6336 10908
rect 6392 10906 6416 10908
rect 6472 10906 6496 10908
rect 6552 10906 6558 10908
rect 6312 10854 6314 10906
rect 6494 10854 6496 10906
rect 6250 10852 6256 10854
rect 6312 10852 6336 10854
rect 6392 10852 6416 10854
rect 6472 10852 6496 10854
rect 6552 10852 6558 10854
rect 6250 10843 6558 10852
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4908 10266 4936 10678
rect 5550 10364 5858 10373
rect 5550 10362 5556 10364
rect 5612 10362 5636 10364
rect 5692 10362 5716 10364
rect 5772 10362 5796 10364
rect 5852 10362 5858 10364
rect 5612 10310 5614 10362
rect 5794 10310 5796 10362
rect 5550 10308 5556 10310
rect 5612 10308 5636 10310
rect 5692 10308 5716 10310
rect 5772 10308 5796 10310
rect 5852 10308 5858 10310
rect 5550 10299 5858 10308
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 6932 10130 6960 11290
rect 7024 11150 7052 11478
rect 7550 11452 7858 11461
rect 7550 11450 7556 11452
rect 7612 11450 7636 11452
rect 7692 11450 7716 11452
rect 7772 11450 7796 11452
rect 7852 11450 7858 11452
rect 7612 11398 7614 11450
rect 7794 11398 7796 11450
rect 7550 11396 7556 11398
rect 7612 11396 7636 11398
rect 7692 11396 7716 11398
rect 7772 11396 7796 11398
rect 7852 11396 7858 11398
rect 7550 11387 7858 11396
rect 8772 11354 8800 11630
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 9232 11218 9260 11630
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4250 9820 4558 9829
rect 4250 9818 4256 9820
rect 4312 9818 4336 9820
rect 4392 9818 4416 9820
rect 4472 9818 4496 9820
rect 4552 9818 4558 9820
rect 4312 9766 4314 9818
rect 4494 9766 4496 9818
rect 4250 9764 4256 9766
rect 4312 9764 4336 9766
rect 4392 9764 4416 9766
rect 4472 9764 4496 9766
rect 4552 9764 4558 9766
rect 4250 9755 4558 9764
rect 4632 9382 4660 9998
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 8906 4660 9318
rect 5356 8968 5408 8974
rect 5460 8945 5488 9590
rect 5550 9276 5858 9285
rect 5550 9274 5556 9276
rect 5612 9274 5636 9276
rect 5692 9274 5716 9276
rect 5772 9274 5796 9276
rect 5852 9274 5858 9276
rect 5612 9222 5614 9274
rect 5794 9222 5796 9274
rect 5550 9220 5556 9222
rect 5612 9220 5636 9222
rect 5692 9220 5716 9222
rect 5772 9220 5796 9222
rect 5852 9220 5858 9222
rect 5550 9211 5858 9220
rect 5920 9178 5948 9930
rect 6250 9820 6558 9829
rect 6250 9818 6256 9820
rect 6312 9818 6336 9820
rect 6392 9818 6416 9820
rect 6472 9818 6496 9820
rect 6552 9818 6558 9820
rect 6312 9766 6314 9818
rect 6494 9766 6496 9818
rect 6250 9764 6256 9766
rect 6312 9764 6336 9766
rect 6392 9764 6416 9766
rect 6472 9764 6496 9766
rect 6552 9764 6558 9766
rect 6250 9755 6558 9764
rect 6932 9674 6960 10066
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6748 9646 6960 9674
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6104 9178 6132 9318
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 5920 9030 6224 9058
rect 5920 8974 5948 9030
rect 5908 8968 5960 8974
rect 5356 8910 5408 8916
rect 5446 8936 5502 8945
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4250 8732 4558 8741
rect 4250 8730 4256 8732
rect 4312 8730 4336 8732
rect 4392 8730 4416 8732
rect 4472 8730 4496 8732
rect 4552 8730 4558 8732
rect 4312 8678 4314 8730
rect 4494 8678 4496 8730
rect 4250 8676 4256 8678
rect 4312 8676 4336 8678
rect 4392 8676 4416 8678
rect 4472 8676 4496 8678
rect 4552 8676 4558 8678
rect 4250 8667 4558 8676
rect 5368 8634 5396 8910
rect 5908 8910 5960 8916
rect 6000 8968 6052 8974
rect 6092 8968 6144 8974
rect 6000 8910 6052 8916
rect 6090 8936 6092 8945
rect 6144 8936 6146 8945
rect 5446 8871 5502 8880
rect 5460 8838 5488 8871
rect 6012 8838 6040 8910
rect 6196 8906 6224 9030
rect 6090 8871 6146 8880
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 6012 8294 6040 8774
rect 6250 8732 6558 8741
rect 6250 8730 6256 8732
rect 6312 8730 6336 8732
rect 6392 8730 6416 8732
rect 6472 8730 6496 8732
rect 6552 8730 6558 8732
rect 6312 8678 6314 8730
rect 6494 8678 6496 8730
rect 6250 8676 6256 8678
rect 6312 8676 6336 8678
rect 6392 8676 6416 8678
rect 6472 8676 6496 8678
rect 6552 8676 6558 8678
rect 6250 8667 6558 8676
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5550 8188 5858 8197
rect 5550 8186 5556 8188
rect 5612 8186 5636 8188
rect 5692 8186 5716 8188
rect 5772 8186 5796 8188
rect 5852 8186 5858 8188
rect 5612 8134 5614 8186
rect 5794 8134 5796 8186
rect 5550 8132 5556 8134
rect 5612 8132 5636 8134
rect 5692 8132 5716 8134
rect 5772 8132 5796 8134
rect 5852 8132 5858 8134
rect 5550 8123 5858 8132
rect 6656 8090 6684 9590
rect 6748 8974 6776 9646
rect 6932 9586 6960 9646
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7024 9518 7052 11086
rect 8250 10908 8558 10917
rect 8250 10906 8256 10908
rect 8312 10906 8336 10908
rect 8392 10906 8416 10908
rect 8472 10906 8496 10908
rect 8552 10906 8558 10908
rect 8312 10854 8314 10906
rect 8494 10854 8496 10906
rect 8250 10852 8256 10854
rect 8312 10852 8336 10854
rect 8392 10852 8416 10854
rect 8472 10852 8496 10854
rect 8552 10852 8558 10854
rect 8250 10843 8558 10852
rect 8588 10554 8616 11154
rect 9324 11098 9352 12174
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9508 11830 9536 12038
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 10060 11762 10088 12038
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9550 11452 9858 11461
rect 9550 11450 9556 11452
rect 9612 11450 9636 11452
rect 9692 11450 9716 11452
rect 9772 11450 9796 11452
rect 9852 11450 9858 11452
rect 9612 11398 9614 11450
rect 9794 11398 9796 11450
rect 9550 11396 9556 11398
rect 9612 11396 9636 11398
rect 9692 11396 9716 11398
rect 9772 11396 9796 11398
rect 9852 11396 9858 11398
rect 9550 11387 9858 11396
rect 9968 11150 9996 11494
rect 10060 11218 10088 11562
rect 10152 11286 10180 12582
rect 10336 12170 10364 12786
rect 10796 12714 10824 12951
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10250 11996 10558 12005
rect 10250 11994 10256 11996
rect 10312 11994 10336 11996
rect 10392 11994 10416 11996
rect 10472 11994 10496 11996
rect 10552 11994 10558 11996
rect 10312 11942 10314 11994
rect 10494 11942 10496 11994
rect 10250 11940 10256 11942
rect 10312 11940 10336 11942
rect 10392 11940 10416 11942
rect 10472 11940 10496 11942
rect 10552 11940 10558 11942
rect 10250 11931 10558 11940
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9232 11070 9352 11098
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8496 10526 8616 10554
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 7550 10364 7858 10373
rect 7550 10362 7556 10364
rect 7612 10362 7636 10364
rect 7692 10362 7716 10364
rect 7772 10362 7796 10364
rect 7852 10362 7858 10364
rect 7612 10310 7614 10362
rect 7794 10310 7796 10362
rect 7550 10308 7556 10310
rect 7612 10308 7636 10310
rect 7692 10308 7716 10310
rect 7772 10308 7796 10310
rect 7852 10308 7858 10310
rect 7550 10299 7858 10308
rect 8496 10062 8524 10526
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8588 10062 8616 10406
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8680 9926 8708 10542
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8498 6776 8910
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 2044 6384 2096 6390
rect 3332 6384 3384 6390
rect 2044 6326 2096 6332
rect 3252 6344 3332 6372
rect 848 6112 900 6118
rect 846 6080 848 6089
rect 900 6080 902 6089
rect 846 6015 902 6024
rect 1550 6012 1858 6021
rect 1550 6010 1556 6012
rect 1612 6010 1636 6012
rect 1692 6010 1716 6012
rect 1772 6010 1796 6012
rect 1852 6010 1858 6012
rect 1612 5958 1614 6010
rect 1794 5958 1796 6010
rect 1550 5956 1556 5958
rect 1612 5956 1636 5958
rect 1692 5956 1716 5958
rect 1772 5956 1796 5958
rect 1852 5956 1858 5958
rect 1550 5947 1858 5956
rect 1964 5914 1992 6326
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2056 5794 2084 6326
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2608 6118 2636 6190
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 1872 5766 2084 5794
rect 848 5568 900 5574
rect 848 5510 900 5516
rect 860 5409 888 5510
rect 846 5400 902 5409
rect 846 5335 902 5344
rect 1872 5166 1900 5766
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1550 4924 1858 4933
rect 1550 4922 1556 4924
rect 1612 4922 1636 4924
rect 1692 4922 1716 4924
rect 1772 4922 1796 4924
rect 1852 4922 1858 4924
rect 1612 4870 1614 4922
rect 1794 4870 1796 4922
rect 1550 4868 1556 4870
rect 1612 4868 1636 4870
rect 1692 4868 1716 4870
rect 1772 4868 1796 4870
rect 1852 4868 1858 4870
rect 1550 4859 1858 4868
rect 1550 3836 1858 3845
rect 1550 3834 1556 3836
rect 1612 3834 1636 3836
rect 1692 3834 1716 3836
rect 1772 3834 1796 3836
rect 1852 3834 1858 3836
rect 1612 3782 1614 3834
rect 1794 3782 1796 3834
rect 1550 3780 1556 3782
rect 1612 3780 1636 3782
rect 1692 3780 1716 3782
rect 1772 3780 1796 3782
rect 1852 3780 1858 3782
rect 1550 3771 1858 3780
rect 1964 3738 1992 5510
rect 2148 5166 2176 5578
rect 2250 5468 2558 5477
rect 2250 5466 2256 5468
rect 2312 5466 2336 5468
rect 2392 5466 2416 5468
rect 2472 5466 2496 5468
rect 2552 5466 2558 5468
rect 2312 5414 2314 5466
rect 2494 5414 2496 5466
rect 2250 5412 2256 5414
rect 2312 5412 2336 5414
rect 2392 5412 2416 5414
rect 2472 5412 2496 5414
rect 2552 5412 2558 5414
rect 2250 5403 2558 5412
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2608 4554 2636 6054
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2884 5778 2912 5850
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2884 5234 2912 5714
rect 2976 5574 3004 6122
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 3068 4826 3096 6122
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5778 3188 6054
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3252 4604 3280 6344
rect 3332 6326 3384 6332
rect 3436 6322 3464 7686
rect 4250 7644 4558 7653
rect 4250 7642 4256 7644
rect 4312 7642 4336 7644
rect 4392 7642 4416 7644
rect 4472 7642 4496 7644
rect 4552 7642 4558 7644
rect 4312 7590 4314 7642
rect 4494 7590 4496 7642
rect 4250 7588 4256 7590
rect 4312 7588 4336 7590
rect 4392 7588 4416 7590
rect 4472 7588 4496 7590
rect 4552 7588 4558 7590
rect 4250 7579 4558 7588
rect 6250 7644 6558 7653
rect 6250 7642 6256 7644
rect 6312 7642 6336 7644
rect 6392 7642 6416 7644
rect 6472 7642 6496 7644
rect 6552 7642 6558 7644
rect 6312 7590 6314 7642
rect 6494 7590 6496 7642
rect 6250 7588 6256 7590
rect 6312 7588 6336 7590
rect 6392 7588 6416 7590
rect 6472 7588 6496 7590
rect 6552 7588 6558 7590
rect 6250 7579 6558 7588
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3550 7100 3858 7109
rect 3550 7098 3556 7100
rect 3612 7098 3636 7100
rect 3692 7098 3716 7100
rect 3772 7098 3796 7100
rect 3852 7098 3858 7100
rect 3612 7046 3614 7098
rect 3794 7046 3796 7098
rect 3550 7044 3556 7046
rect 3612 7044 3636 7046
rect 3692 7044 3716 7046
rect 3772 7044 3796 7046
rect 3852 7044 3858 7046
rect 3550 7035 3858 7044
rect 3988 6322 4016 7346
rect 5550 7100 5858 7109
rect 5550 7098 5556 7100
rect 5612 7098 5636 7100
rect 5692 7098 5716 7100
rect 5772 7098 5796 7100
rect 5852 7098 5858 7100
rect 5612 7046 5614 7098
rect 5794 7046 5796 7098
rect 5550 7044 5556 7046
rect 5612 7044 5636 7046
rect 5692 7044 5716 7046
rect 5772 7044 5796 7046
rect 5852 7044 5858 7046
rect 5550 7035 5858 7044
rect 4250 6556 4558 6565
rect 4250 6554 4256 6556
rect 4312 6554 4336 6556
rect 4392 6554 4416 6556
rect 4472 6554 4496 6556
rect 4552 6554 4558 6556
rect 4312 6502 4314 6554
rect 4494 6502 4496 6554
rect 4250 6500 4256 6502
rect 4312 6500 4336 6502
rect 4392 6500 4416 6502
rect 4472 6500 4496 6502
rect 4552 6500 4558 6502
rect 4250 6491 4558 6500
rect 6250 6556 6558 6565
rect 6250 6554 6256 6556
rect 6312 6554 6336 6556
rect 6392 6554 6416 6556
rect 6472 6554 6496 6556
rect 6552 6554 6558 6556
rect 6312 6502 6314 6554
rect 6494 6502 6496 6554
rect 6250 6500 6256 6502
rect 6312 6500 6336 6502
rect 6392 6500 6416 6502
rect 6472 6500 6496 6502
rect 6552 6500 6558 6502
rect 6250 6491 6558 6500
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3436 6202 3464 6258
rect 3344 6174 3464 6202
rect 3344 5302 3372 6174
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5642 3464 6054
rect 3550 6012 3858 6021
rect 3550 6010 3556 6012
rect 3612 6010 3636 6012
rect 3692 6010 3716 6012
rect 3772 6010 3796 6012
rect 3852 6010 3858 6012
rect 3612 5958 3614 6010
rect 3794 5958 3796 6010
rect 3550 5956 3556 5958
rect 3612 5956 3636 5958
rect 3692 5956 3716 5958
rect 3772 5956 3796 5958
rect 3852 5956 3858 5958
rect 3550 5947 3858 5956
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 5370 3924 5510
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 3344 4758 3372 5238
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 3436 4690 3464 5170
rect 3550 4924 3858 4933
rect 3550 4922 3556 4924
rect 3612 4922 3636 4924
rect 3692 4922 3716 4924
rect 3772 4922 3796 4924
rect 3852 4922 3858 4924
rect 3612 4870 3614 4922
rect 3794 4870 3796 4922
rect 3550 4868 3556 4870
rect 3612 4868 3636 4870
rect 3692 4868 3716 4870
rect 3772 4868 3796 4870
rect 3852 4868 3858 4870
rect 3550 4859 3858 4868
rect 3896 4690 3924 5306
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3332 4616 3384 4622
rect 3252 4576 3332 4604
rect 3988 4570 4016 6258
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5710 4200 6054
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4250 5468 4558 5477
rect 4250 5466 4256 5468
rect 4312 5466 4336 5468
rect 4392 5466 4416 5468
rect 4472 5466 4496 5468
rect 4552 5466 4558 5468
rect 4312 5414 4314 5466
rect 4494 5414 4496 5466
rect 4250 5412 4256 5414
rect 4312 5412 4336 5414
rect 4392 5412 4416 5414
rect 4472 5412 4496 5414
rect 4552 5412 4558 5414
rect 4250 5403 4558 5412
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4080 4622 4108 5306
rect 4908 5234 4936 6326
rect 5092 5370 5120 6326
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 3332 4558 3384 4564
rect 2596 4548 2648 4554
rect 2596 4490 2648 4496
rect 3896 4542 4016 4570
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 2250 4380 2558 4389
rect 2250 4378 2256 4380
rect 2312 4378 2336 4380
rect 2392 4378 2416 4380
rect 2472 4378 2496 4380
rect 2552 4378 2558 4380
rect 2312 4326 2314 4378
rect 2494 4326 2496 4378
rect 2250 4324 2256 4326
rect 2312 4324 2336 4326
rect 2392 4324 2416 4326
rect 2472 4324 2496 4326
rect 2552 4324 2558 4326
rect 2250 4315 2558 4324
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1964 3126 1992 3674
rect 2136 3460 2188 3466
rect 2136 3402 2188 3408
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 2148 2990 2176 3402
rect 2250 3292 2558 3301
rect 2250 3290 2256 3292
rect 2312 3290 2336 3292
rect 2392 3290 2416 3292
rect 2472 3290 2496 3292
rect 2552 3290 2558 3292
rect 2312 3238 2314 3290
rect 2494 3238 2496 3290
rect 2250 3236 2256 3238
rect 2312 3236 2336 3238
rect 2392 3236 2416 3238
rect 2472 3236 2496 3238
rect 2552 3236 2558 3238
rect 2250 3227 2558 3236
rect 2608 2990 2636 4490
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4078 3280 4422
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2700 3194 2728 3878
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 3058 2820 3878
rect 3436 3398 3464 4014
rect 3896 4010 3924 4542
rect 4080 4162 4108 4558
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3988 4134 4108 4162
rect 4172 4146 4200 4422
rect 4250 4380 4558 4389
rect 4250 4378 4256 4380
rect 4312 4378 4336 4380
rect 4392 4378 4416 4380
rect 4472 4378 4496 4380
rect 4552 4378 4558 4380
rect 4312 4326 4314 4378
rect 4494 4326 4496 4378
rect 4250 4324 4256 4326
rect 4312 4324 4336 4326
rect 4392 4324 4416 4326
rect 4472 4324 4496 4326
rect 4552 4324 4558 4326
rect 4250 4315 4558 4324
rect 4160 4140 4212 4146
rect 3988 4078 4016 4134
rect 4160 4082 4212 4088
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3550 3836 3858 3845
rect 3550 3834 3556 3836
rect 3612 3834 3636 3836
rect 3692 3834 3716 3836
rect 3772 3834 3796 3836
rect 3852 3834 3858 3836
rect 3612 3782 3614 3834
rect 3794 3782 3796 3834
rect 3550 3780 3556 3782
rect 3612 3780 3636 3782
rect 3692 3780 3716 3782
rect 3772 3780 3796 3782
rect 3852 3780 3858 3782
rect 3550 3771 3858 3780
rect 4172 3602 4200 4082
rect 4632 4078 4660 5170
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4264 3482 4292 3946
rect 4172 3466 4292 3482
rect 4160 3460 4292 3466
rect 4212 3454 4292 3460
rect 4160 3402 4212 3408
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 1550 2748 1858 2757
rect 1550 2746 1556 2748
rect 1612 2746 1636 2748
rect 1692 2746 1716 2748
rect 1772 2746 1796 2748
rect 1852 2746 1858 2748
rect 1612 2694 1614 2746
rect 1794 2694 1796 2746
rect 1550 2692 1556 2694
rect 1612 2692 1636 2694
rect 1692 2692 1716 2694
rect 1772 2692 1796 2694
rect 1852 2692 1858 2694
rect 1550 2683 1858 2692
rect 3436 2446 3464 3334
rect 3550 2748 3858 2757
rect 3550 2746 3556 2748
rect 3612 2746 3636 2748
rect 3692 2746 3716 2748
rect 3772 2746 3796 2748
rect 3852 2746 3858 2748
rect 3612 2694 3614 2746
rect 3794 2694 3796 2746
rect 3550 2692 3556 2694
rect 3612 2692 3636 2694
rect 3692 2692 3716 2694
rect 3772 2692 3796 2694
rect 3852 2692 3858 2694
rect 3550 2683 3858 2692
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 4172 2378 4200 3402
rect 4250 3292 4558 3301
rect 4250 3290 4256 3292
rect 4312 3290 4336 3292
rect 4392 3290 4416 3292
rect 4472 3290 4496 3292
rect 4552 3290 4558 3292
rect 4312 3238 4314 3290
rect 4494 3238 4496 3290
rect 4250 3236 4256 3238
rect 4312 3236 4336 3238
rect 4392 3236 4416 3238
rect 4472 3236 4496 3238
rect 4552 3236 4558 3238
rect 4250 3227 4558 3236
rect 4632 3194 4660 4014
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5184 3466 5212 3878
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4448 2650 4476 3062
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4632 2514 4660 3130
rect 4724 2990 4752 3402
rect 5368 3194 5396 6054
rect 5550 6012 5858 6021
rect 5550 6010 5556 6012
rect 5612 6010 5636 6012
rect 5692 6010 5716 6012
rect 5772 6010 5796 6012
rect 5852 6010 5858 6012
rect 5612 5958 5614 6010
rect 5794 5958 5796 6010
rect 5550 5956 5556 5958
rect 5612 5956 5636 5958
rect 5692 5956 5716 5958
rect 5772 5956 5796 5958
rect 5852 5956 5858 5958
rect 5550 5947 5858 5956
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 3602 5488 5510
rect 5920 5370 5948 5578
rect 6250 5468 6558 5477
rect 6250 5466 6256 5468
rect 6312 5466 6336 5468
rect 6392 5466 6416 5468
rect 6472 5466 6496 5468
rect 6552 5466 6558 5468
rect 6312 5414 6314 5466
rect 6494 5414 6496 5466
rect 6250 5412 6256 5414
rect 6312 5412 6336 5414
rect 6392 5412 6416 5414
rect 6472 5412 6496 5414
rect 6552 5412 6558 5414
rect 6250 5403 6558 5412
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 5550 4924 5858 4933
rect 5550 4922 5556 4924
rect 5612 4922 5636 4924
rect 5692 4922 5716 4924
rect 5772 4922 5796 4924
rect 5852 4922 5858 4924
rect 5612 4870 5614 4922
rect 5794 4870 5796 4922
rect 5550 4868 5556 4870
rect 5612 4868 5636 4870
rect 5692 4868 5716 4870
rect 5772 4868 5796 4870
rect 5852 4868 5858 4870
rect 5550 4859 5858 4868
rect 5920 4298 5948 5170
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5736 4282 5948 4298
rect 5724 4276 5948 4282
rect 5776 4270 5948 4276
rect 5724 4218 5776 4224
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5550 3836 5858 3845
rect 5550 3834 5556 3836
rect 5612 3834 5636 3836
rect 5692 3834 5716 3836
rect 5772 3834 5796 3836
rect 5852 3834 5858 3836
rect 5612 3782 5614 3834
rect 5794 3782 5796 3834
rect 5550 3780 5556 3782
rect 5612 3780 5636 3782
rect 5692 3780 5716 3782
rect 5772 3780 5796 3782
rect 5852 3780 5858 3782
rect 5550 3771 5858 3780
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5368 2990 5396 3130
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 5356 2984 5408 2990
rect 5828 2972 5856 3334
rect 5920 3126 5948 3878
rect 6012 3738 6040 4626
rect 6656 4554 6684 8026
rect 7024 7886 7052 9454
rect 7300 9042 7328 9862
rect 8128 9704 8156 9862
rect 8250 9820 8558 9829
rect 8250 9818 8256 9820
rect 8312 9818 8336 9820
rect 8392 9818 8416 9820
rect 8472 9818 8496 9820
rect 8552 9818 8558 9820
rect 8312 9766 8314 9818
rect 8494 9766 8496 9818
rect 8250 9764 8256 9766
rect 8312 9764 8336 9766
rect 8392 9764 8416 9766
rect 8472 9764 8496 9766
rect 8552 9764 8558 9766
rect 8250 9755 8558 9764
rect 8128 9676 8248 9704
rect 7654 9616 7710 9625
rect 7654 9551 7656 9560
rect 7708 9551 7710 9560
rect 7656 9522 7708 9528
rect 8220 9518 8248 9676
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7550 9276 7858 9285
rect 7550 9274 7556 9276
rect 7612 9274 7636 9276
rect 7692 9274 7716 9276
rect 7772 9274 7796 9276
rect 7852 9274 7858 9276
rect 7612 9222 7614 9274
rect 7794 9222 7796 9274
rect 7550 9220 7556 9222
rect 7612 9220 7636 9222
rect 7692 9220 7716 9222
rect 7772 9220 7796 9222
rect 7852 9220 7858 9222
rect 7550 9211 7858 9220
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7944 8906 7972 9318
rect 8680 9178 8708 9862
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 8024 8832 8076 8838
rect 7944 8780 8024 8786
rect 7944 8774 8076 8780
rect 7944 8758 8064 8774
rect 7944 8498 7972 8758
rect 8250 8732 8558 8741
rect 8250 8730 8256 8732
rect 8312 8730 8336 8732
rect 8392 8730 8416 8732
rect 8472 8730 8496 8732
rect 8552 8730 8558 8732
rect 8312 8678 8314 8730
rect 8494 8678 8496 8730
rect 8250 8676 8256 8678
rect 8312 8676 8336 8678
rect 8392 8676 8416 8678
rect 8472 8676 8496 8678
rect 8552 8676 8558 8678
rect 8250 8667 8558 8676
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 7954 7328 8230
rect 7550 8188 7858 8197
rect 7550 8186 7556 8188
rect 7612 8186 7636 8188
rect 7692 8186 7716 8188
rect 7772 8186 7796 8188
rect 7852 8186 7858 8188
rect 7612 8134 7614 8186
rect 7794 8134 7796 8186
rect 7550 8132 7556 8134
rect 7612 8132 7636 8134
rect 7692 8132 7716 8134
rect 7772 8132 7796 8134
rect 7852 8132 7858 8134
rect 7550 8123 7858 8132
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 7410 7052 7822
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7300 7002 7328 7278
rect 7550 7100 7858 7109
rect 7550 7098 7556 7100
rect 7612 7098 7636 7100
rect 7692 7098 7716 7100
rect 7772 7098 7796 7100
rect 7852 7098 7858 7100
rect 7612 7046 7614 7098
rect 7794 7046 7796 7098
rect 7550 7044 7556 7046
rect 7612 7044 7636 7046
rect 7692 7044 7716 7046
rect 7772 7044 7796 7046
rect 7852 7044 7858 7046
rect 7550 7035 7858 7044
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7944 6866 7972 8434
rect 8250 7644 8558 7653
rect 8250 7642 8256 7644
rect 8312 7642 8336 7644
rect 8392 7642 8416 7644
rect 8472 7642 8496 7644
rect 8552 7642 8558 7644
rect 8312 7590 8314 7642
rect 8494 7590 8496 7642
rect 8250 7588 8256 7590
rect 8312 7588 8336 7590
rect 8392 7588 8416 7590
rect 8472 7588 8496 7590
rect 8552 7588 8558 7590
rect 8250 7579 8558 7588
rect 8680 7546 8708 8570
rect 8772 8566 8800 10610
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 8772 7886 8800 8502
rect 8864 8090 8892 10066
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 8956 9722 8984 9930
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 9048 9625 9076 10610
rect 9034 9616 9090 9625
rect 9034 9551 9090 9560
rect 9048 8906 9076 9551
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9036 8424 9088 8430
rect 9034 8392 9036 8401
rect 9088 8392 9090 8401
rect 9034 8327 9090 8336
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 9048 8022 9076 8327
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9140 7886 9168 8774
rect 9232 8498 9260 11070
rect 9968 10742 9996 11086
rect 10250 10908 10558 10917
rect 10250 10906 10256 10908
rect 10312 10906 10336 10908
rect 10392 10906 10416 10908
rect 10472 10906 10496 10908
rect 10552 10906 10558 10908
rect 10312 10854 10314 10906
rect 10494 10854 10496 10906
rect 10250 10852 10256 10854
rect 10312 10852 10336 10854
rect 10392 10852 10416 10854
rect 10472 10852 10496 10854
rect 10552 10852 10558 10854
rect 10250 10843 10558 10852
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 9586 9352 10406
rect 9550 10364 9858 10373
rect 9550 10362 9556 10364
rect 9612 10362 9636 10364
rect 9692 10362 9716 10364
rect 9772 10362 9796 10364
rect 9852 10362 9858 10364
rect 9612 10310 9614 10362
rect 9794 10310 9796 10362
rect 9550 10308 9556 10310
rect 9612 10308 9636 10310
rect 9692 10308 9716 10310
rect 9772 10308 9796 10310
rect 9852 10308 9858 10310
rect 9550 10299 9858 10308
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9784 9654 9812 9998
rect 9968 9926 9996 10678
rect 10612 10606 10640 12310
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10704 11694 10732 12106
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9232 8022 9260 8434
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9416 7970 9444 9386
rect 9550 9276 9858 9285
rect 9550 9274 9556 9276
rect 9612 9274 9636 9276
rect 9692 9274 9716 9276
rect 9772 9274 9796 9276
rect 9852 9274 9858 9276
rect 9612 9222 9614 9274
rect 9794 9222 9796 9274
rect 9550 9220 9556 9222
rect 9612 9220 9636 9222
rect 9692 9220 9716 9222
rect 9772 9220 9796 9222
rect 9852 9220 9858 9222
rect 9550 9211 9858 9220
rect 9968 9042 9996 9862
rect 10250 9820 10558 9829
rect 10250 9818 10256 9820
rect 10312 9818 10336 9820
rect 10392 9818 10416 9820
rect 10472 9818 10496 9820
rect 10552 9818 10558 9820
rect 10312 9766 10314 9818
rect 10494 9766 10496 9818
rect 10250 9764 10256 9766
rect 10312 9764 10336 9766
rect 10392 9764 10416 9766
rect 10472 9764 10496 9766
rect 10552 9764 10558 9766
rect 10250 9755 10558 9764
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10060 9178 10088 9590
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9508 8430 9536 8842
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9600 8498 9628 8570
rect 9876 8566 9904 8774
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9586 8392 9642 8401
rect 9586 8327 9588 8336
rect 9640 8327 9642 8336
rect 9588 8298 9640 8304
rect 9550 8188 9858 8197
rect 9550 8186 9556 8188
rect 9612 8186 9636 8188
rect 9692 8186 9716 8188
rect 9772 8186 9796 8188
rect 9852 8186 9858 8188
rect 9612 8134 9614 8186
rect 9794 8134 9796 8186
rect 9550 8132 9556 8134
rect 9612 8132 9636 8134
rect 9692 8132 9716 8134
rect 9772 8132 9796 8134
rect 9852 8132 9858 8134
rect 9550 8123 9858 8132
rect 9968 8090 9996 8842
rect 10060 8634 10088 8910
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10250 8732 10558 8741
rect 10250 8730 10256 8732
rect 10312 8730 10336 8732
rect 10392 8730 10416 8732
rect 10472 8730 10496 8732
rect 10552 8730 10558 8732
rect 10312 8678 10314 8730
rect 10494 8678 10496 8730
rect 10250 8676 10256 8678
rect 10312 8676 10336 8678
rect 10392 8676 10416 8678
rect 10472 8676 10496 8678
rect 10552 8676 10558 8678
rect 10250 8667 10558 8676
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10140 8560 10192 8566
rect 10138 8528 10140 8537
rect 10192 8528 10194 8537
rect 10704 8498 10732 8774
rect 10796 8634 10824 9862
rect 10888 9654 10916 11698
rect 10980 10062 11008 11766
rect 11072 11082 11100 12854
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 12345 11192 12582
rect 11150 12336 11206 12345
rect 11150 12271 11206 12280
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11164 10742 11192 11698
rect 11256 11626 11284 12786
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11348 11830 11376 12582
rect 11550 12540 11858 12549
rect 11550 12538 11556 12540
rect 11612 12538 11636 12540
rect 11692 12538 11716 12540
rect 11772 12538 11796 12540
rect 11852 12538 11858 12540
rect 11612 12486 11614 12538
rect 11794 12486 11796 12538
rect 11550 12484 11556 12486
rect 11612 12484 11636 12486
rect 11692 12484 11716 12486
rect 11772 12484 11796 12486
rect 11852 12484 11858 12486
rect 11550 12475 11858 12484
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11440 10810 11468 12174
rect 11992 11665 12020 12582
rect 12084 12442 12112 12786
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 11978 11656 12034 11665
rect 11978 11591 12034 11600
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11550 11452 11858 11461
rect 11550 11450 11556 11452
rect 11612 11450 11636 11452
rect 11692 11450 11716 11452
rect 11772 11450 11796 11452
rect 11852 11450 11858 11452
rect 11612 11398 11614 11450
rect 11794 11398 11796 11450
rect 11550 11396 11556 11398
rect 11612 11396 11636 11398
rect 11692 11396 11716 11398
rect 11772 11396 11796 11398
rect 11852 11396 11858 11398
rect 11550 11387 11858 11396
rect 11900 10985 11928 11494
rect 12084 11354 12112 12378
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11886 10976 11942 10985
rect 11886 10911 11942 10920
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10980 9586 11008 9998
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10138 8463 10194 8472
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9416 7942 9536 7970
rect 9508 7886 9536 7942
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8680 7410 8708 7482
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 6932 5302 6960 6802
rect 8312 6798 8340 7210
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8250 6556 8558 6565
rect 8250 6554 8256 6556
rect 8312 6554 8336 6556
rect 8392 6554 8416 6556
rect 8472 6554 8496 6556
rect 8552 6554 8558 6556
rect 8312 6502 8314 6554
rect 8494 6502 8496 6554
rect 8250 6500 8256 6502
rect 8312 6500 8336 6502
rect 8392 6500 8416 6502
rect 8472 6500 8496 6502
rect 8552 6500 8558 6502
rect 8250 6491 8558 6500
rect 8864 6458 8892 6734
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 7550 6012 7858 6021
rect 7550 6010 7556 6012
rect 7612 6010 7636 6012
rect 7692 6010 7716 6012
rect 7772 6010 7796 6012
rect 7852 6010 7858 6012
rect 7612 5958 7614 6010
rect 7794 5958 7796 6010
rect 7550 5956 7556 5958
rect 7612 5956 7636 5958
rect 7692 5956 7716 5958
rect 7772 5956 7796 5958
rect 7852 5956 7858 5958
rect 7550 5947 7858 5956
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7300 5574 7328 5646
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6250 4380 6558 4389
rect 6250 4378 6256 4380
rect 6312 4378 6336 4380
rect 6392 4378 6416 4380
rect 6472 4378 6496 4380
rect 6552 4378 6558 4380
rect 6312 4326 6314 4378
rect 6494 4326 6496 4378
rect 6250 4324 6256 4326
rect 6312 4324 6336 4326
rect 6392 4324 6416 4326
rect 6472 4324 6496 4326
rect 6552 4324 6558 4326
rect 6250 4315 6558 4324
rect 6092 4208 6144 4214
rect 6144 4156 6316 4162
rect 6092 4150 6316 4156
rect 6104 4134 6316 4150
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6012 3126 6040 3674
rect 6196 3482 6224 3946
rect 6288 3602 6316 4134
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6196 3466 6408 3482
rect 6184 3460 6408 3466
rect 6236 3454 6408 3460
rect 6184 3402 6236 3408
rect 6380 3398 6408 3454
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5828 2944 5948 2972
rect 5356 2926 5408 2932
rect 5920 2774 5948 2944
rect 6104 2854 6132 3334
rect 6250 3292 6558 3301
rect 6250 3290 6256 3292
rect 6312 3290 6336 3292
rect 6392 3290 6416 3292
rect 6472 3290 6496 3292
rect 6552 3290 6558 3292
rect 6312 3238 6314 3290
rect 6494 3238 6496 3290
rect 6250 3236 6256 3238
rect 6312 3236 6336 3238
rect 6392 3236 6416 3238
rect 6472 3236 6496 3238
rect 6552 3236 6558 3238
rect 6250 3227 6558 3236
rect 6748 3058 6776 3538
rect 6840 3194 6868 5170
rect 7116 4690 7144 5170
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7300 4282 7328 5510
rect 7484 5302 7512 5510
rect 8128 5302 8156 5578
rect 8250 5468 8558 5477
rect 8250 5466 8256 5468
rect 8312 5466 8336 5468
rect 8392 5466 8416 5468
rect 8472 5466 8496 5468
rect 8552 5466 8558 5468
rect 8312 5414 8314 5466
rect 8494 5414 8496 5466
rect 8250 5412 8256 5414
rect 8312 5412 8336 5414
rect 8392 5412 8416 5414
rect 8472 5412 8496 5414
rect 8552 5412 8558 5414
rect 8250 5403 8558 5412
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 7550 4924 7858 4933
rect 7550 4922 7556 4924
rect 7612 4922 7636 4924
rect 7692 4922 7716 4924
rect 7772 4922 7796 4924
rect 7852 4922 7858 4924
rect 7612 4870 7614 4922
rect 7794 4870 7796 4922
rect 7550 4868 7556 4870
rect 7612 4868 7636 4870
rect 7692 4868 7716 4870
rect 7772 4868 7796 4870
rect 7852 4868 7858 4870
rect 7550 4859 7858 4868
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6380 2854 6408 2926
rect 6092 2848 6144 2854
rect 6092 2790 6144 2796
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 5550 2748 5858 2757
rect 5550 2746 5556 2748
rect 5612 2746 5636 2748
rect 5692 2746 5716 2748
rect 5772 2746 5796 2748
rect 5852 2746 5858 2748
rect 5920 2746 6040 2774
rect 5612 2694 5614 2746
rect 5794 2694 5796 2746
rect 5550 2692 5556 2694
rect 5612 2692 5636 2694
rect 5692 2692 5716 2694
rect 5772 2692 5796 2694
rect 5852 2692 5858 2694
rect 5550 2683 5858 2692
rect 6012 2514 6040 2746
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6748 2446 6776 2994
rect 6932 2854 6960 4150
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 2582 6960 2790
rect 7024 2650 7052 2858
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 7116 2446 7144 3062
rect 7300 2446 7328 4218
rect 7392 4146 7420 4762
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8036 4146 8064 4626
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7550 3836 7858 3845
rect 7550 3834 7556 3836
rect 7612 3834 7636 3836
rect 7692 3834 7716 3836
rect 7772 3834 7796 3836
rect 7852 3834 7858 3836
rect 7612 3782 7614 3834
rect 7794 3782 7796 3834
rect 7550 3780 7556 3782
rect 7612 3780 7636 3782
rect 7692 3780 7716 3782
rect 7772 3780 7796 3782
rect 7852 3780 7858 3782
rect 7550 3771 7858 3780
rect 8128 3738 8156 4558
rect 8250 4380 8558 4389
rect 8250 4378 8256 4380
rect 8312 4378 8336 4380
rect 8392 4378 8416 4380
rect 8472 4378 8496 4380
rect 8552 4378 8558 4380
rect 8312 4326 8314 4378
rect 8494 4326 8496 4378
rect 8250 4324 8256 4326
rect 8312 4324 8336 4326
rect 8392 4324 8416 4326
rect 8472 4324 8496 4326
rect 8552 4324 8558 4326
rect 8250 4315 8558 4324
rect 8588 4162 8616 5714
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5302 8708 5510
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8956 5166 8984 6802
rect 9048 5778 9076 7278
rect 9550 7100 9858 7109
rect 9550 7098 9556 7100
rect 9612 7098 9636 7100
rect 9692 7098 9716 7100
rect 9772 7098 9796 7100
rect 9852 7098 9858 7100
rect 9612 7046 9614 7098
rect 9794 7046 9796 7098
rect 9550 7044 9556 7046
rect 9612 7044 9636 7046
rect 9692 7044 9716 7046
rect 9772 7044 9796 7046
rect 9852 7044 9858 7046
rect 9550 7035 9858 7044
rect 9968 6934 9996 7890
rect 10060 7886 10088 8366
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 7954 10364 8230
rect 10888 8090 10916 8842
rect 11072 8090 11100 10542
rect 11440 10062 11468 10746
rect 12084 10538 12112 11290
rect 12176 10810 12204 12038
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 11550 10364 11858 10373
rect 11550 10362 11556 10364
rect 11612 10362 11636 10364
rect 11692 10362 11716 10364
rect 11772 10362 11796 10364
rect 11852 10362 11858 10364
rect 11612 10310 11614 10362
rect 11794 10310 11796 10362
rect 11550 10308 11556 10310
rect 11612 10308 11636 10310
rect 11692 10308 11716 10310
rect 11772 10308 11796 10310
rect 11852 10308 11858 10310
rect 11550 10299 11858 10308
rect 11978 10296 12034 10305
rect 11978 10231 11980 10240
rect 12032 10231 12034 10240
rect 11980 10202 12032 10208
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11164 8838 11192 9454
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11164 8566 11192 8774
rect 11256 8634 11284 9930
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11152 8560 11204 8566
rect 11348 8537 11376 9930
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11152 8502 11204 8508
rect 11334 8528 11390 8537
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11164 8022 11192 8502
rect 11440 8498 11468 9862
rect 12070 9616 12126 9625
rect 12176 9586 12204 10746
rect 12070 9551 12126 9560
rect 12164 9580 12216 9586
rect 11550 9276 11858 9285
rect 11550 9274 11556 9276
rect 11612 9274 11636 9276
rect 11692 9274 11716 9276
rect 11772 9274 11796 9276
rect 11852 9274 11858 9276
rect 11612 9222 11614 9274
rect 11794 9222 11796 9274
rect 11550 9220 11556 9222
rect 11612 9220 11636 9222
rect 11692 9220 11716 9222
rect 11772 9220 11796 9222
rect 11852 9220 11858 9222
rect 11550 9211 11858 9220
rect 11886 8936 11942 8945
rect 11886 8871 11942 8880
rect 11334 8463 11390 8472
rect 11428 8492 11480 8498
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 11348 7886 11376 8463
rect 11428 8434 11480 8440
rect 11550 8188 11858 8197
rect 11550 8186 11556 8188
rect 11612 8186 11636 8188
rect 11692 8186 11716 8188
rect 11772 8186 11796 8188
rect 11852 8186 11858 8188
rect 11612 8134 11614 8186
rect 11794 8134 11796 8186
rect 11550 8132 11556 8134
rect 11612 8132 11636 8134
rect 11692 8132 11716 8134
rect 11772 8132 11796 8134
rect 11852 8132 11858 8134
rect 11550 8123 11858 8132
rect 11900 8090 11928 8871
rect 12084 8634 12112 9551
rect 12164 9522 12216 9528
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12176 8430 12204 9522
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 12084 8265 12112 8298
rect 12070 8256 12126 8265
rect 12070 8191 12126 8200
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 10250 7644 10558 7653
rect 10250 7642 10256 7644
rect 10312 7642 10336 7644
rect 10392 7642 10416 7644
rect 10472 7642 10496 7644
rect 10552 7642 10558 7644
rect 10312 7590 10314 7642
rect 10494 7590 10496 7642
rect 10250 7588 10256 7590
rect 10312 7588 10336 7590
rect 10392 7588 10416 7590
rect 10472 7588 10496 7590
rect 10552 7588 10558 7590
rect 10250 7579 10558 7588
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9968 6390 9996 6734
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9416 5386 9444 6190
rect 9550 6012 9858 6021
rect 9550 6010 9556 6012
rect 9612 6010 9636 6012
rect 9692 6010 9716 6012
rect 9772 6010 9796 6012
rect 9852 6010 9858 6012
rect 9612 5958 9614 6010
rect 9794 5958 9796 6010
rect 9550 5956 9556 5958
rect 9612 5956 9636 5958
rect 9692 5956 9716 5958
rect 9772 5956 9796 5958
rect 9852 5956 9858 5958
rect 9550 5947 9858 5956
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9416 5370 9536 5386
rect 9416 5364 9548 5370
rect 9416 5358 9496 5364
rect 9496 5306 9548 5312
rect 9784 5234 9812 5782
rect 9968 5642 9996 6326
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5914 10088 6054
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 9550 4924 9858 4933
rect 9550 4922 9556 4924
rect 9612 4922 9636 4924
rect 9692 4922 9716 4924
rect 9772 4922 9796 4924
rect 9852 4922 9858 4924
rect 9612 4870 9614 4922
rect 9794 4870 9796 4922
rect 9550 4868 9556 4870
rect 9612 4868 9636 4870
rect 9692 4868 9716 4870
rect 9772 4868 9796 4870
rect 9852 4868 9858 4870
rect 9550 4859 9858 4868
rect 9968 4826 9996 5578
rect 10152 5370 10180 6666
rect 10250 6556 10558 6565
rect 10250 6554 10256 6556
rect 10312 6554 10336 6556
rect 10392 6554 10416 6556
rect 10472 6554 10496 6556
rect 10552 6554 10558 6556
rect 10312 6502 10314 6554
rect 10494 6502 10496 6554
rect 10250 6500 10256 6502
rect 10312 6500 10336 6502
rect 10392 6500 10416 6502
rect 10472 6500 10496 6502
rect 10552 6500 10558 6502
rect 10250 6491 10558 6500
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10250 5468 10558 5477
rect 10250 5466 10256 5468
rect 10312 5466 10336 5468
rect 10392 5466 10416 5468
rect 10472 5466 10496 5468
rect 10552 5466 10558 5468
rect 10312 5414 10314 5466
rect 10494 5414 10496 5466
rect 10250 5412 10256 5414
rect 10312 5412 10336 5414
rect 10392 5412 10416 5414
rect 10472 5412 10496 5414
rect 10552 5412 10558 5414
rect 10250 5403 10558 5412
rect 10612 5370 10640 6326
rect 10796 5778 10824 6802
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9404 4548 9456 4554
rect 9404 4490 9456 4496
rect 9416 4282 9444 4490
rect 9508 4282 9536 4694
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 8496 4134 8616 4162
rect 9508 4146 9536 4218
rect 9496 4140 9548 4146
rect 8496 4078 8524 4134
rect 9496 4082 9548 4088
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8496 3534 8524 4014
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 7392 2650 7420 3470
rect 7656 3392 7708 3398
rect 7576 3340 7656 3346
rect 7576 3334 7708 3340
rect 7576 3318 7696 3334
rect 7576 3126 7604 3318
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7550 2748 7858 2757
rect 7550 2746 7556 2748
rect 7612 2746 7636 2748
rect 7692 2746 7716 2748
rect 7772 2746 7796 2748
rect 7852 2746 7858 2748
rect 7612 2694 7614 2746
rect 7794 2694 7796 2746
rect 7550 2692 7556 2694
rect 7612 2692 7636 2694
rect 7692 2692 7716 2694
rect 7772 2692 7796 2694
rect 7852 2692 7858 2694
rect 7550 2683 7858 2692
rect 7944 2650 7972 2926
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8036 2446 8064 3470
rect 8250 3292 8558 3301
rect 8250 3290 8256 3292
rect 8312 3290 8336 3292
rect 8392 3290 8416 3292
rect 8472 3290 8496 3292
rect 8552 3290 8558 3292
rect 8312 3238 8314 3290
rect 8494 3238 8496 3290
rect 8250 3236 8256 3238
rect 8312 3236 8336 3238
rect 8392 3236 8416 3238
rect 8472 3236 8496 3238
rect 8552 3236 8558 3238
rect 8250 3227 8558 3236
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9048 2650 9076 2994
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9232 2514 9260 3878
rect 9416 3534 9444 3878
rect 9550 3836 9858 3845
rect 9550 3834 9556 3836
rect 9612 3834 9636 3836
rect 9692 3834 9716 3836
rect 9772 3834 9796 3836
rect 9852 3834 9858 3836
rect 9612 3782 9614 3834
rect 9794 3782 9796 3834
rect 9550 3780 9556 3782
rect 9612 3780 9636 3782
rect 9692 3780 9716 3782
rect 9772 3780 9796 3782
rect 9852 3780 9858 3782
rect 9550 3771 9858 3780
rect 9968 3602 9996 4762
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9876 2990 9904 3402
rect 9968 3126 9996 3538
rect 10060 3466 10088 4966
rect 10152 4078 10180 5170
rect 10244 4486 10272 5170
rect 10704 5098 10732 5714
rect 10796 5302 10824 5714
rect 10980 5642 11008 7346
rect 11164 6186 11192 7822
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11440 7585 11468 7686
rect 11426 7576 11482 7585
rect 11426 7511 11482 7520
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11256 6730 11284 7142
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11256 5778 11284 6054
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10980 5522 11008 5578
rect 10980 5494 11100 5522
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10796 4826 10824 5238
rect 11072 5234 11100 5494
rect 11256 5370 11284 5714
rect 11348 5642 11376 7142
rect 11550 7100 11858 7109
rect 11550 7098 11556 7100
rect 11612 7098 11636 7100
rect 11692 7098 11716 7100
rect 11772 7098 11796 7100
rect 11852 7098 11858 7100
rect 11612 7046 11614 7098
rect 11794 7046 11796 7098
rect 11550 7044 11556 7046
rect 11612 7044 11636 7046
rect 11692 7044 11716 7046
rect 11772 7044 11796 7046
rect 11852 7044 11858 7046
rect 11550 7035 11858 7044
rect 11900 6905 11928 7142
rect 11886 6896 11942 6905
rect 11886 6831 11942 6840
rect 11992 6662 12020 7278
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11072 5030 11100 5170
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10250 4380 10558 4389
rect 10250 4378 10256 4380
rect 10312 4378 10336 4380
rect 10392 4378 10416 4380
rect 10472 4378 10496 4380
rect 10552 4378 10558 4380
rect 10312 4326 10314 4378
rect 10494 4326 10496 4378
rect 10250 4324 10256 4326
rect 10312 4324 10336 4326
rect 10392 4324 10416 4326
rect 10472 4324 10496 4326
rect 10552 4324 10558 4326
rect 10250 4315 10558 4324
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10428 4078 10456 4218
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3602 10456 4014
rect 10704 3738 10732 4422
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10250 3292 10558 3301
rect 10250 3290 10256 3292
rect 10312 3290 10336 3292
rect 10392 3290 10416 3292
rect 10472 3290 10496 3292
rect 10552 3290 10558 3292
rect 10312 3238 10314 3290
rect 10494 3238 10496 3290
rect 10250 3236 10256 3238
rect 10312 3236 10336 3238
rect 10392 3236 10416 3238
rect 10472 3236 10496 3238
rect 10552 3236 10558 3238
rect 10250 3227 10558 3236
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9550 2748 9858 2757
rect 9550 2746 9556 2748
rect 9612 2746 9636 2748
rect 9692 2746 9716 2748
rect 9772 2746 9796 2748
rect 9852 2746 9858 2748
rect 9612 2694 9614 2746
rect 9794 2694 9796 2746
rect 9550 2692 9556 2694
rect 9612 2692 9636 2694
rect 9692 2692 9716 2694
rect 9772 2692 9796 2694
rect 9852 2692 9858 2694
rect 9550 2683 9858 2692
rect 9968 2514 9996 2790
rect 10704 2650 10732 3402
rect 10980 2922 11008 3538
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 11072 2446 11100 4966
rect 11164 4690 11192 5238
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11256 4622 11284 5306
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11164 4146 11192 4490
rect 11348 4486 11376 4966
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11164 3738 11192 4082
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11440 3194 11468 6258
rect 11886 6216 11942 6225
rect 11886 6151 11942 6160
rect 11550 6012 11858 6021
rect 11550 6010 11556 6012
rect 11612 6010 11636 6012
rect 11692 6010 11716 6012
rect 11772 6010 11796 6012
rect 11852 6010 11858 6012
rect 11612 5958 11614 6010
rect 11794 5958 11796 6010
rect 11550 5956 11556 5958
rect 11612 5956 11636 5958
rect 11692 5956 11716 5958
rect 11772 5956 11796 5958
rect 11852 5956 11858 5958
rect 11550 5947 11858 5956
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5302 11836 5510
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11550 4924 11858 4933
rect 11550 4922 11556 4924
rect 11612 4922 11636 4924
rect 11692 4922 11716 4924
rect 11772 4922 11796 4924
rect 11852 4922 11858 4924
rect 11612 4870 11614 4922
rect 11794 4870 11796 4922
rect 11550 4868 11556 4870
rect 11612 4868 11636 4870
rect 11692 4868 11716 4870
rect 11772 4868 11796 4870
rect 11852 4868 11858 4870
rect 11550 4859 11858 4868
rect 11900 4826 11928 6151
rect 11992 5098 12020 6598
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12070 5536 12126 5545
rect 12070 5471 12126 5480
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 11978 4856 12034 4865
rect 11888 4820 11940 4826
rect 11978 4791 12034 4800
rect 11888 4762 11940 4768
rect 11794 4176 11850 4185
rect 11794 4111 11850 4120
rect 11808 4010 11836 4111
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 11550 3836 11858 3845
rect 11550 3834 11556 3836
rect 11612 3834 11636 3836
rect 11692 3834 11716 3836
rect 11772 3834 11796 3836
rect 11852 3834 11858 3836
rect 11612 3782 11614 3834
rect 11794 3782 11796 3834
rect 11550 3780 11556 3782
rect 11612 3780 11636 3782
rect 11692 3780 11716 3782
rect 11772 3780 11796 3782
rect 11852 3780 11858 3782
rect 11550 3771 11858 3780
rect 11794 3496 11850 3505
rect 11794 3431 11850 3440
rect 11808 3398 11836 3431
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11256 2650 11284 3062
rect 11992 3058 12020 4791
rect 12084 4758 12112 5471
rect 12176 5234 12204 6054
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12176 4078 12204 5170
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11978 2816 12034 2825
rect 11550 2748 11858 2757
rect 11978 2751 12034 2760
rect 11550 2746 11556 2748
rect 11612 2746 11636 2748
rect 11692 2746 11716 2748
rect 11772 2746 11796 2748
rect 11852 2746 11858 2748
rect 11612 2694 11614 2746
rect 11794 2694 11796 2746
rect 11550 2692 11556 2694
rect 11612 2692 11636 2694
rect 11692 2692 11716 2694
rect 11772 2692 11796 2694
rect 11852 2692 11858 2694
rect 11550 2683 11858 2692
rect 11992 2650 12020 2751
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 2250 2204 2558 2213
rect 2250 2202 2256 2204
rect 2312 2202 2336 2204
rect 2392 2202 2416 2204
rect 2472 2202 2496 2204
rect 2552 2202 2558 2204
rect 2312 2150 2314 2202
rect 2494 2150 2496 2202
rect 2250 2148 2256 2150
rect 2312 2148 2336 2150
rect 2392 2148 2416 2150
rect 2472 2148 2496 2150
rect 2552 2148 2558 2150
rect 2250 2139 2558 2148
rect 3252 800 3280 2246
rect 3896 800 3924 2246
rect 4250 2204 4558 2213
rect 4250 2202 4256 2204
rect 4312 2202 4336 2204
rect 4392 2202 4416 2204
rect 4472 2202 4496 2204
rect 4552 2202 4558 2204
rect 4312 2150 4314 2202
rect 4494 2150 4496 2202
rect 4250 2148 4256 2150
rect 4312 2148 4336 2150
rect 4392 2148 4416 2150
rect 4472 2148 4496 2150
rect 4552 2148 4558 2150
rect 4250 2139 4558 2148
rect 5828 800 5856 2246
rect 6250 2204 6558 2213
rect 6250 2202 6256 2204
rect 6312 2202 6336 2204
rect 6392 2202 6416 2204
rect 6472 2202 6496 2204
rect 6552 2202 6558 2204
rect 6312 2150 6314 2202
rect 6494 2150 6496 2202
rect 6250 2148 6256 2150
rect 6312 2148 6336 2150
rect 6392 2148 6416 2150
rect 6472 2148 6496 2150
rect 6552 2148 6558 2150
rect 6250 2139 6558 2148
rect 6656 1170 6684 2246
rect 6472 1142 6684 1170
rect 6472 800 6500 1142
rect 7116 800 7144 2246
rect 7760 800 7788 2246
rect 8250 2204 8558 2213
rect 8250 2202 8256 2204
rect 8312 2202 8336 2204
rect 8392 2202 8416 2204
rect 8472 2202 8496 2204
rect 8552 2202 8558 2204
rect 8312 2150 8314 2202
rect 8494 2150 8496 2202
rect 8250 2148 8256 2150
rect 8312 2148 8336 2150
rect 8392 2148 8416 2150
rect 8472 2148 8496 2150
rect 8552 2148 8558 2150
rect 8250 2139 8558 2148
rect 9048 800 9076 2246
rect 10250 2204 10558 2213
rect 10250 2202 10256 2204
rect 10312 2202 10336 2204
rect 10392 2202 10416 2204
rect 10472 2202 10496 2204
rect 10552 2202 10558 2204
rect 10312 2150 10314 2202
rect 10494 2150 10496 2202
rect 10250 2148 10256 2150
rect 10312 2148 10336 2150
rect 10392 2148 10416 2150
rect 10472 2148 10496 2150
rect 10552 2148 10558 2150
rect 10250 2139 10558 2148
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 9034 0 9090 800
<< via2 >>
rect 2256 13082 2312 13084
rect 2336 13082 2392 13084
rect 2416 13082 2472 13084
rect 2496 13082 2552 13084
rect 2256 13030 2302 13082
rect 2302 13030 2312 13082
rect 2336 13030 2366 13082
rect 2366 13030 2378 13082
rect 2378 13030 2392 13082
rect 2416 13030 2430 13082
rect 2430 13030 2442 13082
rect 2442 13030 2472 13082
rect 2496 13030 2506 13082
rect 2506 13030 2552 13082
rect 2256 13028 2312 13030
rect 2336 13028 2392 13030
rect 2416 13028 2472 13030
rect 2496 13028 2552 13030
rect 4256 13082 4312 13084
rect 4336 13082 4392 13084
rect 4416 13082 4472 13084
rect 4496 13082 4552 13084
rect 4256 13030 4302 13082
rect 4302 13030 4312 13082
rect 4336 13030 4366 13082
rect 4366 13030 4378 13082
rect 4378 13030 4392 13082
rect 4416 13030 4430 13082
rect 4430 13030 4442 13082
rect 4442 13030 4472 13082
rect 4496 13030 4506 13082
rect 4506 13030 4552 13082
rect 4256 13028 4312 13030
rect 4336 13028 4392 13030
rect 4416 13028 4472 13030
rect 4496 13028 4552 13030
rect 6256 13082 6312 13084
rect 6336 13082 6392 13084
rect 6416 13082 6472 13084
rect 6496 13082 6552 13084
rect 6256 13030 6302 13082
rect 6302 13030 6312 13082
rect 6336 13030 6366 13082
rect 6366 13030 6378 13082
rect 6378 13030 6392 13082
rect 6416 13030 6430 13082
rect 6430 13030 6442 13082
rect 6442 13030 6472 13082
rect 6496 13030 6506 13082
rect 6506 13030 6552 13082
rect 6256 13028 6312 13030
rect 6336 13028 6392 13030
rect 6416 13028 6472 13030
rect 6496 13028 6552 13030
rect 8256 13082 8312 13084
rect 8336 13082 8392 13084
rect 8416 13082 8472 13084
rect 8496 13082 8552 13084
rect 8256 13030 8302 13082
rect 8302 13030 8312 13082
rect 8336 13030 8366 13082
rect 8366 13030 8378 13082
rect 8378 13030 8392 13082
rect 8416 13030 8430 13082
rect 8430 13030 8442 13082
rect 8442 13030 8472 13082
rect 8496 13030 8506 13082
rect 8506 13030 8552 13082
rect 8256 13028 8312 13030
rect 8336 13028 8392 13030
rect 8416 13028 8472 13030
rect 8496 13028 8552 13030
rect 10256 13082 10312 13084
rect 10336 13082 10392 13084
rect 10416 13082 10472 13084
rect 10496 13082 10552 13084
rect 10256 13030 10302 13082
rect 10302 13030 10312 13082
rect 10336 13030 10366 13082
rect 10366 13030 10378 13082
rect 10378 13030 10392 13082
rect 10416 13030 10430 13082
rect 10430 13030 10442 13082
rect 10442 13030 10472 13082
rect 10496 13030 10506 13082
rect 10506 13030 10552 13082
rect 10256 13028 10312 13030
rect 10336 13028 10392 13030
rect 10416 13028 10472 13030
rect 10496 13028 10552 13030
rect 10782 12960 10838 13016
rect 1556 12538 1612 12540
rect 1636 12538 1692 12540
rect 1716 12538 1772 12540
rect 1796 12538 1852 12540
rect 1556 12486 1602 12538
rect 1602 12486 1612 12538
rect 1636 12486 1666 12538
rect 1666 12486 1678 12538
rect 1678 12486 1692 12538
rect 1716 12486 1730 12538
rect 1730 12486 1742 12538
rect 1742 12486 1772 12538
rect 1796 12486 1806 12538
rect 1806 12486 1852 12538
rect 1556 12484 1612 12486
rect 1636 12484 1692 12486
rect 1716 12484 1772 12486
rect 1796 12484 1852 12486
rect 3556 12538 3612 12540
rect 3636 12538 3692 12540
rect 3716 12538 3772 12540
rect 3796 12538 3852 12540
rect 3556 12486 3602 12538
rect 3602 12486 3612 12538
rect 3636 12486 3666 12538
rect 3666 12486 3678 12538
rect 3678 12486 3692 12538
rect 3716 12486 3730 12538
rect 3730 12486 3742 12538
rect 3742 12486 3772 12538
rect 3796 12486 3806 12538
rect 3806 12486 3852 12538
rect 3556 12484 3612 12486
rect 3636 12484 3692 12486
rect 3716 12484 3772 12486
rect 3796 12484 3852 12486
rect 2256 11994 2312 11996
rect 2336 11994 2392 11996
rect 2416 11994 2472 11996
rect 2496 11994 2552 11996
rect 2256 11942 2302 11994
rect 2302 11942 2312 11994
rect 2336 11942 2366 11994
rect 2366 11942 2378 11994
rect 2378 11942 2392 11994
rect 2416 11942 2430 11994
rect 2430 11942 2442 11994
rect 2442 11942 2472 11994
rect 2496 11942 2506 11994
rect 2506 11942 2552 11994
rect 2256 11940 2312 11942
rect 2336 11940 2392 11942
rect 2416 11940 2472 11942
rect 2496 11940 2552 11942
rect 1556 11450 1612 11452
rect 1636 11450 1692 11452
rect 1716 11450 1772 11452
rect 1796 11450 1852 11452
rect 1556 11398 1602 11450
rect 1602 11398 1612 11450
rect 1636 11398 1666 11450
rect 1666 11398 1678 11450
rect 1678 11398 1692 11450
rect 1716 11398 1730 11450
rect 1730 11398 1742 11450
rect 1742 11398 1772 11450
rect 1796 11398 1806 11450
rect 1806 11398 1852 11450
rect 1556 11396 1612 11398
rect 1636 11396 1692 11398
rect 1716 11396 1772 11398
rect 1796 11396 1852 11398
rect 1556 10362 1612 10364
rect 1636 10362 1692 10364
rect 1716 10362 1772 10364
rect 1796 10362 1852 10364
rect 1556 10310 1602 10362
rect 1602 10310 1612 10362
rect 1636 10310 1666 10362
rect 1666 10310 1678 10362
rect 1678 10310 1692 10362
rect 1716 10310 1730 10362
rect 1730 10310 1742 10362
rect 1742 10310 1772 10362
rect 1796 10310 1806 10362
rect 1806 10310 1852 10362
rect 1556 10308 1612 10310
rect 1636 10308 1692 10310
rect 1716 10308 1772 10310
rect 1796 10308 1852 10310
rect 2256 10906 2312 10908
rect 2336 10906 2392 10908
rect 2416 10906 2472 10908
rect 2496 10906 2552 10908
rect 2256 10854 2302 10906
rect 2302 10854 2312 10906
rect 2336 10854 2366 10906
rect 2366 10854 2378 10906
rect 2378 10854 2392 10906
rect 2416 10854 2430 10906
rect 2430 10854 2442 10906
rect 2442 10854 2472 10906
rect 2496 10854 2506 10906
rect 2506 10854 2552 10906
rect 2256 10852 2312 10854
rect 2336 10852 2392 10854
rect 2416 10852 2472 10854
rect 2496 10852 2552 10854
rect 3556 11450 3612 11452
rect 3636 11450 3692 11452
rect 3716 11450 3772 11452
rect 3796 11450 3852 11452
rect 3556 11398 3602 11450
rect 3602 11398 3612 11450
rect 3636 11398 3666 11450
rect 3666 11398 3678 11450
rect 3678 11398 3692 11450
rect 3716 11398 3730 11450
rect 3730 11398 3742 11450
rect 3742 11398 3772 11450
rect 3796 11398 3806 11450
rect 3806 11398 3852 11450
rect 3556 11396 3612 11398
rect 3636 11396 3692 11398
rect 3716 11396 3772 11398
rect 3796 11396 3852 11398
rect 3556 10362 3612 10364
rect 3636 10362 3692 10364
rect 3716 10362 3772 10364
rect 3796 10362 3852 10364
rect 3556 10310 3602 10362
rect 3602 10310 3612 10362
rect 3636 10310 3666 10362
rect 3666 10310 3678 10362
rect 3678 10310 3692 10362
rect 3716 10310 3730 10362
rect 3730 10310 3742 10362
rect 3742 10310 3772 10362
rect 3796 10310 3806 10362
rect 3806 10310 3852 10362
rect 3556 10308 3612 10310
rect 3636 10308 3692 10310
rect 3716 10308 3772 10310
rect 3796 10308 3852 10310
rect 846 9424 902 9480
rect 846 9052 848 9072
rect 848 9052 900 9072
rect 900 9052 902 9072
rect 846 9016 902 9052
rect 1556 9274 1612 9276
rect 1636 9274 1692 9276
rect 1716 9274 1772 9276
rect 1796 9274 1852 9276
rect 1556 9222 1602 9274
rect 1602 9222 1612 9274
rect 1636 9222 1666 9274
rect 1666 9222 1678 9274
rect 1678 9222 1692 9274
rect 1716 9222 1730 9274
rect 1730 9222 1742 9274
rect 1742 9222 1772 9274
rect 1796 9222 1806 9274
rect 1806 9222 1852 9274
rect 1556 9220 1612 9222
rect 1636 9220 1692 9222
rect 1716 9220 1772 9222
rect 1796 9220 1852 9222
rect 846 8064 902 8120
rect 846 7692 848 7712
rect 848 7692 900 7712
rect 900 7692 902 7712
rect 846 7656 902 7692
rect 2256 9818 2312 9820
rect 2336 9818 2392 9820
rect 2416 9818 2472 9820
rect 2496 9818 2552 9820
rect 2256 9766 2302 9818
rect 2302 9766 2312 9818
rect 2336 9766 2366 9818
rect 2366 9766 2378 9818
rect 2378 9766 2392 9818
rect 2416 9766 2430 9818
rect 2430 9766 2442 9818
rect 2442 9766 2472 9818
rect 2496 9766 2506 9818
rect 2506 9766 2552 9818
rect 2256 9764 2312 9766
rect 2336 9764 2392 9766
rect 2416 9764 2472 9766
rect 2496 9764 2552 9766
rect 4256 11994 4312 11996
rect 4336 11994 4392 11996
rect 4416 11994 4472 11996
rect 4496 11994 4552 11996
rect 4256 11942 4302 11994
rect 4302 11942 4312 11994
rect 4336 11942 4366 11994
rect 4366 11942 4378 11994
rect 4378 11942 4392 11994
rect 4416 11942 4430 11994
rect 4430 11942 4442 11994
rect 4442 11942 4472 11994
rect 4496 11942 4506 11994
rect 4506 11942 4552 11994
rect 4256 11940 4312 11942
rect 4336 11940 4392 11942
rect 4416 11940 4472 11942
rect 4496 11940 4552 11942
rect 4158 11600 4214 11656
rect 5556 12538 5612 12540
rect 5636 12538 5692 12540
rect 5716 12538 5772 12540
rect 5796 12538 5852 12540
rect 5556 12486 5602 12538
rect 5602 12486 5612 12538
rect 5636 12486 5666 12538
rect 5666 12486 5678 12538
rect 5678 12486 5692 12538
rect 5716 12486 5730 12538
rect 5730 12486 5742 12538
rect 5742 12486 5772 12538
rect 5796 12486 5806 12538
rect 5806 12486 5852 12538
rect 5556 12484 5612 12486
rect 5636 12484 5692 12486
rect 5716 12484 5772 12486
rect 5796 12484 5852 12486
rect 2256 8730 2312 8732
rect 2336 8730 2392 8732
rect 2416 8730 2472 8732
rect 2496 8730 2552 8732
rect 2256 8678 2302 8730
rect 2302 8678 2312 8730
rect 2336 8678 2366 8730
rect 2366 8678 2378 8730
rect 2378 8678 2392 8730
rect 2416 8678 2430 8730
rect 2430 8678 2442 8730
rect 2442 8678 2472 8730
rect 2496 8678 2506 8730
rect 2506 8678 2552 8730
rect 2256 8676 2312 8678
rect 2336 8676 2392 8678
rect 2416 8676 2472 8678
rect 2496 8676 2552 8678
rect 1556 8186 1612 8188
rect 1636 8186 1692 8188
rect 1716 8186 1772 8188
rect 1796 8186 1852 8188
rect 1556 8134 1602 8186
rect 1602 8134 1612 8186
rect 1636 8134 1666 8186
rect 1666 8134 1678 8186
rect 1678 8134 1692 8186
rect 1716 8134 1730 8186
rect 1730 8134 1742 8186
rect 1742 8134 1772 8186
rect 1796 8134 1806 8186
rect 1806 8134 1852 8186
rect 1556 8132 1612 8134
rect 1636 8132 1692 8134
rect 1716 8132 1772 8134
rect 1796 8132 1852 8134
rect 3556 9274 3612 9276
rect 3636 9274 3692 9276
rect 3716 9274 3772 9276
rect 3796 9274 3852 9276
rect 3556 9222 3602 9274
rect 3602 9222 3612 9274
rect 3636 9222 3666 9274
rect 3666 9222 3678 9274
rect 3678 9222 3692 9274
rect 3716 9222 3730 9274
rect 3730 9222 3742 9274
rect 3742 9222 3772 9274
rect 3796 9222 3806 9274
rect 3806 9222 3852 9274
rect 3556 9220 3612 9222
rect 3636 9220 3692 9222
rect 3716 9220 3772 9222
rect 3796 9220 3852 9222
rect 2256 7642 2312 7644
rect 2336 7642 2392 7644
rect 2416 7642 2472 7644
rect 2496 7642 2552 7644
rect 2256 7590 2302 7642
rect 2302 7590 2312 7642
rect 2336 7590 2366 7642
rect 2366 7590 2378 7642
rect 2378 7590 2392 7642
rect 2416 7590 2430 7642
rect 2430 7590 2442 7642
rect 2442 7590 2472 7642
rect 2496 7590 2506 7642
rect 2506 7590 2552 7642
rect 2256 7588 2312 7590
rect 2336 7588 2392 7590
rect 2416 7588 2472 7590
rect 2496 7588 2552 7590
rect 1556 7098 1612 7100
rect 1636 7098 1692 7100
rect 1716 7098 1772 7100
rect 1796 7098 1852 7100
rect 1556 7046 1602 7098
rect 1602 7046 1612 7098
rect 1636 7046 1666 7098
rect 1666 7046 1678 7098
rect 1678 7046 1692 7098
rect 1716 7046 1730 7098
rect 1730 7046 1742 7098
rect 1742 7046 1772 7098
rect 1796 7046 1806 7098
rect 1806 7046 1852 7098
rect 1556 7044 1612 7046
rect 1636 7044 1692 7046
rect 1716 7044 1772 7046
rect 1796 7044 1852 7046
rect 2256 6554 2312 6556
rect 2336 6554 2392 6556
rect 2416 6554 2472 6556
rect 2496 6554 2552 6556
rect 2256 6502 2302 6554
rect 2302 6502 2312 6554
rect 2336 6502 2366 6554
rect 2366 6502 2378 6554
rect 2378 6502 2392 6554
rect 2416 6502 2430 6554
rect 2430 6502 2442 6554
rect 2442 6502 2472 6554
rect 2496 6502 2506 6554
rect 2506 6502 2552 6554
rect 2256 6500 2312 6502
rect 2336 6500 2392 6502
rect 2416 6500 2472 6502
rect 2496 6500 2552 6502
rect 3556 8186 3612 8188
rect 3636 8186 3692 8188
rect 3716 8186 3772 8188
rect 3796 8186 3852 8188
rect 3556 8134 3602 8186
rect 3602 8134 3612 8186
rect 3636 8134 3666 8186
rect 3666 8134 3678 8186
rect 3678 8134 3692 8186
rect 3716 8134 3730 8186
rect 3730 8134 3742 8186
rect 3742 8134 3772 8186
rect 3796 8134 3806 8186
rect 3806 8134 3852 8186
rect 3556 8132 3612 8134
rect 3636 8132 3692 8134
rect 3716 8132 3772 8134
rect 3796 8132 3852 8134
rect 4256 10906 4312 10908
rect 4336 10906 4392 10908
rect 4416 10906 4472 10908
rect 4496 10906 4552 10908
rect 4256 10854 4302 10906
rect 4302 10854 4312 10906
rect 4336 10854 4366 10906
rect 4366 10854 4378 10906
rect 4378 10854 4392 10906
rect 4416 10854 4430 10906
rect 4430 10854 4442 10906
rect 4442 10854 4472 10906
rect 4496 10854 4506 10906
rect 4506 10854 4552 10906
rect 4256 10852 4312 10854
rect 4336 10852 4392 10854
rect 4416 10852 4472 10854
rect 4496 10852 4552 10854
rect 6256 11994 6312 11996
rect 6336 11994 6392 11996
rect 6416 11994 6472 11996
rect 6496 11994 6552 11996
rect 6256 11942 6302 11994
rect 6302 11942 6312 11994
rect 6336 11942 6366 11994
rect 6366 11942 6378 11994
rect 6378 11942 6392 11994
rect 6416 11942 6430 11994
rect 6430 11942 6442 11994
rect 6442 11942 6472 11994
rect 6496 11942 6506 11994
rect 6506 11942 6552 11994
rect 6256 11940 6312 11942
rect 6336 11940 6392 11942
rect 6416 11940 6472 11942
rect 6496 11940 6552 11942
rect 5556 11450 5612 11452
rect 5636 11450 5692 11452
rect 5716 11450 5772 11452
rect 5796 11450 5852 11452
rect 5556 11398 5602 11450
rect 5602 11398 5612 11450
rect 5636 11398 5666 11450
rect 5666 11398 5678 11450
rect 5678 11398 5692 11450
rect 5716 11398 5730 11450
rect 5730 11398 5742 11450
rect 5742 11398 5772 11450
rect 5796 11398 5806 11450
rect 5806 11398 5852 11450
rect 5556 11396 5612 11398
rect 5636 11396 5692 11398
rect 5716 11396 5772 11398
rect 5796 11396 5852 11398
rect 7556 12538 7612 12540
rect 7636 12538 7692 12540
rect 7716 12538 7772 12540
rect 7796 12538 7852 12540
rect 7556 12486 7602 12538
rect 7602 12486 7612 12538
rect 7636 12486 7666 12538
rect 7666 12486 7678 12538
rect 7678 12486 7692 12538
rect 7716 12486 7730 12538
rect 7730 12486 7742 12538
rect 7742 12486 7772 12538
rect 7796 12486 7806 12538
rect 7806 12486 7852 12538
rect 7556 12484 7612 12486
rect 7636 12484 7692 12486
rect 7716 12484 7772 12486
rect 7796 12484 7852 12486
rect 9556 12538 9612 12540
rect 9636 12538 9692 12540
rect 9716 12538 9772 12540
rect 9796 12538 9852 12540
rect 9556 12486 9602 12538
rect 9602 12486 9612 12538
rect 9636 12486 9666 12538
rect 9666 12486 9678 12538
rect 9678 12486 9692 12538
rect 9716 12486 9730 12538
rect 9730 12486 9742 12538
rect 9742 12486 9772 12538
rect 9796 12486 9806 12538
rect 9806 12486 9852 12538
rect 9556 12484 9612 12486
rect 9636 12484 9692 12486
rect 9716 12484 9772 12486
rect 9796 12484 9852 12486
rect 8256 11994 8312 11996
rect 8336 11994 8392 11996
rect 8416 11994 8472 11996
rect 8496 11994 8552 11996
rect 8256 11942 8302 11994
rect 8302 11942 8312 11994
rect 8336 11942 8366 11994
rect 8366 11942 8378 11994
rect 8378 11942 8392 11994
rect 8416 11942 8430 11994
rect 8430 11942 8442 11994
rect 8442 11942 8472 11994
rect 8496 11942 8506 11994
rect 8506 11942 8552 11994
rect 8256 11940 8312 11942
rect 8336 11940 8392 11942
rect 8416 11940 8472 11942
rect 8496 11940 8552 11942
rect 6256 10906 6312 10908
rect 6336 10906 6392 10908
rect 6416 10906 6472 10908
rect 6496 10906 6552 10908
rect 6256 10854 6302 10906
rect 6302 10854 6312 10906
rect 6336 10854 6366 10906
rect 6366 10854 6378 10906
rect 6378 10854 6392 10906
rect 6416 10854 6430 10906
rect 6430 10854 6442 10906
rect 6442 10854 6472 10906
rect 6496 10854 6506 10906
rect 6506 10854 6552 10906
rect 6256 10852 6312 10854
rect 6336 10852 6392 10854
rect 6416 10852 6472 10854
rect 6496 10852 6552 10854
rect 5556 10362 5612 10364
rect 5636 10362 5692 10364
rect 5716 10362 5772 10364
rect 5796 10362 5852 10364
rect 5556 10310 5602 10362
rect 5602 10310 5612 10362
rect 5636 10310 5666 10362
rect 5666 10310 5678 10362
rect 5678 10310 5692 10362
rect 5716 10310 5730 10362
rect 5730 10310 5742 10362
rect 5742 10310 5772 10362
rect 5796 10310 5806 10362
rect 5806 10310 5852 10362
rect 5556 10308 5612 10310
rect 5636 10308 5692 10310
rect 5716 10308 5772 10310
rect 5796 10308 5852 10310
rect 7556 11450 7612 11452
rect 7636 11450 7692 11452
rect 7716 11450 7772 11452
rect 7796 11450 7852 11452
rect 7556 11398 7602 11450
rect 7602 11398 7612 11450
rect 7636 11398 7666 11450
rect 7666 11398 7678 11450
rect 7678 11398 7692 11450
rect 7716 11398 7730 11450
rect 7730 11398 7742 11450
rect 7742 11398 7772 11450
rect 7796 11398 7806 11450
rect 7806 11398 7852 11450
rect 7556 11396 7612 11398
rect 7636 11396 7692 11398
rect 7716 11396 7772 11398
rect 7796 11396 7852 11398
rect 4256 9818 4312 9820
rect 4336 9818 4392 9820
rect 4416 9818 4472 9820
rect 4496 9818 4552 9820
rect 4256 9766 4302 9818
rect 4302 9766 4312 9818
rect 4336 9766 4366 9818
rect 4366 9766 4378 9818
rect 4378 9766 4392 9818
rect 4416 9766 4430 9818
rect 4430 9766 4442 9818
rect 4442 9766 4472 9818
rect 4496 9766 4506 9818
rect 4506 9766 4552 9818
rect 4256 9764 4312 9766
rect 4336 9764 4392 9766
rect 4416 9764 4472 9766
rect 4496 9764 4552 9766
rect 5556 9274 5612 9276
rect 5636 9274 5692 9276
rect 5716 9274 5772 9276
rect 5796 9274 5852 9276
rect 5556 9222 5602 9274
rect 5602 9222 5612 9274
rect 5636 9222 5666 9274
rect 5666 9222 5678 9274
rect 5678 9222 5692 9274
rect 5716 9222 5730 9274
rect 5730 9222 5742 9274
rect 5742 9222 5772 9274
rect 5796 9222 5806 9274
rect 5806 9222 5852 9274
rect 5556 9220 5612 9222
rect 5636 9220 5692 9222
rect 5716 9220 5772 9222
rect 5796 9220 5852 9222
rect 6256 9818 6312 9820
rect 6336 9818 6392 9820
rect 6416 9818 6472 9820
rect 6496 9818 6552 9820
rect 6256 9766 6302 9818
rect 6302 9766 6312 9818
rect 6336 9766 6366 9818
rect 6366 9766 6378 9818
rect 6378 9766 6392 9818
rect 6416 9766 6430 9818
rect 6430 9766 6442 9818
rect 6442 9766 6472 9818
rect 6496 9766 6506 9818
rect 6506 9766 6552 9818
rect 6256 9764 6312 9766
rect 6336 9764 6392 9766
rect 6416 9764 6472 9766
rect 6496 9764 6552 9766
rect 4256 8730 4312 8732
rect 4336 8730 4392 8732
rect 4416 8730 4472 8732
rect 4496 8730 4552 8732
rect 4256 8678 4302 8730
rect 4302 8678 4312 8730
rect 4336 8678 4366 8730
rect 4366 8678 4378 8730
rect 4378 8678 4392 8730
rect 4416 8678 4430 8730
rect 4430 8678 4442 8730
rect 4442 8678 4472 8730
rect 4496 8678 4506 8730
rect 4506 8678 4552 8730
rect 4256 8676 4312 8678
rect 4336 8676 4392 8678
rect 4416 8676 4472 8678
rect 4496 8676 4552 8678
rect 5446 8880 5502 8936
rect 6090 8916 6092 8936
rect 6092 8916 6144 8936
rect 6144 8916 6146 8936
rect 6090 8880 6146 8916
rect 6256 8730 6312 8732
rect 6336 8730 6392 8732
rect 6416 8730 6472 8732
rect 6496 8730 6552 8732
rect 6256 8678 6302 8730
rect 6302 8678 6312 8730
rect 6336 8678 6366 8730
rect 6366 8678 6378 8730
rect 6378 8678 6392 8730
rect 6416 8678 6430 8730
rect 6430 8678 6442 8730
rect 6442 8678 6472 8730
rect 6496 8678 6506 8730
rect 6506 8678 6552 8730
rect 6256 8676 6312 8678
rect 6336 8676 6392 8678
rect 6416 8676 6472 8678
rect 6496 8676 6552 8678
rect 5556 8186 5612 8188
rect 5636 8186 5692 8188
rect 5716 8186 5772 8188
rect 5796 8186 5852 8188
rect 5556 8134 5602 8186
rect 5602 8134 5612 8186
rect 5636 8134 5666 8186
rect 5666 8134 5678 8186
rect 5678 8134 5692 8186
rect 5716 8134 5730 8186
rect 5730 8134 5742 8186
rect 5742 8134 5772 8186
rect 5796 8134 5806 8186
rect 5806 8134 5852 8186
rect 5556 8132 5612 8134
rect 5636 8132 5692 8134
rect 5716 8132 5772 8134
rect 5796 8132 5852 8134
rect 8256 10906 8312 10908
rect 8336 10906 8392 10908
rect 8416 10906 8472 10908
rect 8496 10906 8552 10908
rect 8256 10854 8302 10906
rect 8302 10854 8312 10906
rect 8336 10854 8366 10906
rect 8366 10854 8378 10906
rect 8378 10854 8392 10906
rect 8416 10854 8430 10906
rect 8430 10854 8442 10906
rect 8442 10854 8472 10906
rect 8496 10854 8506 10906
rect 8506 10854 8552 10906
rect 8256 10852 8312 10854
rect 8336 10852 8392 10854
rect 8416 10852 8472 10854
rect 8496 10852 8552 10854
rect 9556 11450 9612 11452
rect 9636 11450 9692 11452
rect 9716 11450 9772 11452
rect 9796 11450 9852 11452
rect 9556 11398 9602 11450
rect 9602 11398 9612 11450
rect 9636 11398 9666 11450
rect 9666 11398 9678 11450
rect 9678 11398 9692 11450
rect 9716 11398 9730 11450
rect 9730 11398 9742 11450
rect 9742 11398 9772 11450
rect 9796 11398 9806 11450
rect 9806 11398 9852 11450
rect 9556 11396 9612 11398
rect 9636 11396 9692 11398
rect 9716 11396 9772 11398
rect 9796 11396 9852 11398
rect 10256 11994 10312 11996
rect 10336 11994 10392 11996
rect 10416 11994 10472 11996
rect 10496 11994 10552 11996
rect 10256 11942 10302 11994
rect 10302 11942 10312 11994
rect 10336 11942 10366 11994
rect 10366 11942 10378 11994
rect 10378 11942 10392 11994
rect 10416 11942 10430 11994
rect 10430 11942 10442 11994
rect 10442 11942 10472 11994
rect 10496 11942 10506 11994
rect 10506 11942 10552 11994
rect 10256 11940 10312 11942
rect 10336 11940 10392 11942
rect 10416 11940 10472 11942
rect 10496 11940 10552 11942
rect 7556 10362 7612 10364
rect 7636 10362 7692 10364
rect 7716 10362 7772 10364
rect 7796 10362 7852 10364
rect 7556 10310 7602 10362
rect 7602 10310 7612 10362
rect 7636 10310 7666 10362
rect 7666 10310 7678 10362
rect 7678 10310 7692 10362
rect 7716 10310 7730 10362
rect 7730 10310 7742 10362
rect 7742 10310 7772 10362
rect 7796 10310 7806 10362
rect 7806 10310 7852 10362
rect 7556 10308 7612 10310
rect 7636 10308 7692 10310
rect 7716 10308 7772 10310
rect 7796 10308 7852 10310
rect 846 6060 848 6080
rect 848 6060 900 6080
rect 900 6060 902 6080
rect 846 6024 902 6060
rect 1556 6010 1612 6012
rect 1636 6010 1692 6012
rect 1716 6010 1772 6012
rect 1796 6010 1852 6012
rect 1556 5958 1602 6010
rect 1602 5958 1612 6010
rect 1636 5958 1666 6010
rect 1666 5958 1678 6010
rect 1678 5958 1692 6010
rect 1716 5958 1730 6010
rect 1730 5958 1742 6010
rect 1742 5958 1772 6010
rect 1796 5958 1806 6010
rect 1806 5958 1852 6010
rect 1556 5956 1612 5958
rect 1636 5956 1692 5958
rect 1716 5956 1772 5958
rect 1796 5956 1852 5958
rect 846 5344 902 5400
rect 1556 4922 1612 4924
rect 1636 4922 1692 4924
rect 1716 4922 1772 4924
rect 1796 4922 1852 4924
rect 1556 4870 1602 4922
rect 1602 4870 1612 4922
rect 1636 4870 1666 4922
rect 1666 4870 1678 4922
rect 1678 4870 1692 4922
rect 1716 4870 1730 4922
rect 1730 4870 1742 4922
rect 1742 4870 1772 4922
rect 1796 4870 1806 4922
rect 1806 4870 1852 4922
rect 1556 4868 1612 4870
rect 1636 4868 1692 4870
rect 1716 4868 1772 4870
rect 1796 4868 1852 4870
rect 1556 3834 1612 3836
rect 1636 3834 1692 3836
rect 1716 3834 1772 3836
rect 1796 3834 1852 3836
rect 1556 3782 1602 3834
rect 1602 3782 1612 3834
rect 1636 3782 1666 3834
rect 1666 3782 1678 3834
rect 1678 3782 1692 3834
rect 1716 3782 1730 3834
rect 1730 3782 1742 3834
rect 1742 3782 1772 3834
rect 1796 3782 1806 3834
rect 1806 3782 1852 3834
rect 1556 3780 1612 3782
rect 1636 3780 1692 3782
rect 1716 3780 1772 3782
rect 1796 3780 1852 3782
rect 2256 5466 2312 5468
rect 2336 5466 2392 5468
rect 2416 5466 2472 5468
rect 2496 5466 2552 5468
rect 2256 5414 2302 5466
rect 2302 5414 2312 5466
rect 2336 5414 2366 5466
rect 2366 5414 2378 5466
rect 2378 5414 2392 5466
rect 2416 5414 2430 5466
rect 2430 5414 2442 5466
rect 2442 5414 2472 5466
rect 2496 5414 2506 5466
rect 2506 5414 2552 5466
rect 2256 5412 2312 5414
rect 2336 5412 2392 5414
rect 2416 5412 2472 5414
rect 2496 5412 2552 5414
rect 4256 7642 4312 7644
rect 4336 7642 4392 7644
rect 4416 7642 4472 7644
rect 4496 7642 4552 7644
rect 4256 7590 4302 7642
rect 4302 7590 4312 7642
rect 4336 7590 4366 7642
rect 4366 7590 4378 7642
rect 4378 7590 4392 7642
rect 4416 7590 4430 7642
rect 4430 7590 4442 7642
rect 4442 7590 4472 7642
rect 4496 7590 4506 7642
rect 4506 7590 4552 7642
rect 4256 7588 4312 7590
rect 4336 7588 4392 7590
rect 4416 7588 4472 7590
rect 4496 7588 4552 7590
rect 6256 7642 6312 7644
rect 6336 7642 6392 7644
rect 6416 7642 6472 7644
rect 6496 7642 6552 7644
rect 6256 7590 6302 7642
rect 6302 7590 6312 7642
rect 6336 7590 6366 7642
rect 6366 7590 6378 7642
rect 6378 7590 6392 7642
rect 6416 7590 6430 7642
rect 6430 7590 6442 7642
rect 6442 7590 6472 7642
rect 6496 7590 6506 7642
rect 6506 7590 6552 7642
rect 6256 7588 6312 7590
rect 6336 7588 6392 7590
rect 6416 7588 6472 7590
rect 6496 7588 6552 7590
rect 3556 7098 3612 7100
rect 3636 7098 3692 7100
rect 3716 7098 3772 7100
rect 3796 7098 3852 7100
rect 3556 7046 3602 7098
rect 3602 7046 3612 7098
rect 3636 7046 3666 7098
rect 3666 7046 3678 7098
rect 3678 7046 3692 7098
rect 3716 7046 3730 7098
rect 3730 7046 3742 7098
rect 3742 7046 3772 7098
rect 3796 7046 3806 7098
rect 3806 7046 3852 7098
rect 3556 7044 3612 7046
rect 3636 7044 3692 7046
rect 3716 7044 3772 7046
rect 3796 7044 3852 7046
rect 5556 7098 5612 7100
rect 5636 7098 5692 7100
rect 5716 7098 5772 7100
rect 5796 7098 5852 7100
rect 5556 7046 5602 7098
rect 5602 7046 5612 7098
rect 5636 7046 5666 7098
rect 5666 7046 5678 7098
rect 5678 7046 5692 7098
rect 5716 7046 5730 7098
rect 5730 7046 5742 7098
rect 5742 7046 5772 7098
rect 5796 7046 5806 7098
rect 5806 7046 5852 7098
rect 5556 7044 5612 7046
rect 5636 7044 5692 7046
rect 5716 7044 5772 7046
rect 5796 7044 5852 7046
rect 4256 6554 4312 6556
rect 4336 6554 4392 6556
rect 4416 6554 4472 6556
rect 4496 6554 4552 6556
rect 4256 6502 4302 6554
rect 4302 6502 4312 6554
rect 4336 6502 4366 6554
rect 4366 6502 4378 6554
rect 4378 6502 4392 6554
rect 4416 6502 4430 6554
rect 4430 6502 4442 6554
rect 4442 6502 4472 6554
rect 4496 6502 4506 6554
rect 4506 6502 4552 6554
rect 4256 6500 4312 6502
rect 4336 6500 4392 6502
rect 4416 6500 4472 6502
rect 4496 6500 4552 6502
rect 6256 6554 6312 6556
rect 6336 6554 6392 6556
rect 6416 6554 6472 6556
rect 6496 6554 6552 6556
rect 6256 6502 6302 6554
rect 6302 6502 6312 6554
rect 6336 6502 6366 6554
rect 6366 6502 6378 6554
rect 6378 6502 6392 6554
rect 6416 6502 6430 6554
rect 6430 6502 6442 6554
rect 6442 6502 6472 6554
rect 6496 6502 6506 6554
rect 6506 6502 6552 6554
rect 6256 6500 6312 6502
rect 6336 6500 6392 6502
rect 6416 6500 6472 6502
rect 6496 6500 6552 6502
rect 3556 6010 3612 6012
rect 3636 6010 3692 6012
rect 3716 6010 3772 6012
rect 3796 6010 3852 6012
rect 3556 5958 3602 6010
rect 3602 5958 3612 6010
rect 3636 5958 3666 6010
rect 3666 5958 3678 6010
rect 3678 5958 3692 6010
rect 3716 5958 3730 6010
rect 3730 5958 3742 6010
rect 3742 5958 3772 6010
rect 3796 5958 3806 6010
rect 3806 5958 3852 6010
rect 3556 5956 3612 5958
rect 3636 5956 3692 5958
rect 3716 5956 3772 5958
rect 3796 5956 3852 5958
rect 3556 4922 3612 4924
rect 3636 4922 3692 4924
rect 3716 4922 3772 4924
rect 3796 4922 3852 4924
rect 3556 4870 3602 4922
rect 3602 4870 3612 4922
rect 3636 4870 3666 4922
rect 3666 4870 3678 4922
rect 3678 4870 3692 4922
rect 3716 4870 3730 4922
rect 3730 4870 3742 4922
rect 3742 4870 3772 4922
rect 3796 4870 3806 4922
rect 3806 4870 3852 4922
rect 3556 4868 3612 4870
rect 3636 4868 3692 4870
rect 3716 4868 3772 4870
rect 3796 4868 3852 4870
rect 4256 5466 4312 5468
rect 4336 5466 4392 5468
rect 4416 5466 4472 5468
rect 4496 5466 4552 5468
rect 4256 5414 4302 5466
rect 4302 5414 4312 5466
rect 4336 5414 4366 5466
rect 4366 5414 4378 5466
rect 4378 5414 4392 5466
rect 4416 5414 4430 5466
rect 4430 5414 4442 5466
rect 4442 5414 4472 5466
rect 4496 5414 4506 5466
rect 4506 5414 4552 5466
rect 4256 5412 4312 5414
rect 4336 5412 4392 5414
rect 4416 5412 4472 5414
rect 4496 5412 4552 5414
rect 2256 4378 2312 4380
rect 2336 4378 2392 4380
rect 2416 4378 2472 4380
rect 2496 4378 2552 4380
rect 2256 4326 2302 4378
rect 2302 4326 2312 4378
rect 2336 4326 2366 4378
rect 2366 4326 2378 4378
rect 2378 4326 2392 4378
rect 2416 4326 2430 4378
rect 2430 4326 2442 4378
rect 2442 4326 2472 4378
rect 2496 4326 2506 4378
rect 2506 4326 2552 4378
rect 2256 4324 2312 4326
rect 2336 4324 2392 4326
rect 2416 4324 2472 4326
rect 2496 4324 2552 4326
rect 2256 3290 2312 3292
rect 2336 3290 2392 3292
rect 2416 3290 2472 3292
rect 2496 3290 2552 3292
rect 2256 3238 2302 3290
rect 2302 3238 2312 3290
rect 2336 3238 2366 3290
rect 2366 3238 2378 3290
rect 2378 3238 2392 3290
rect 2416 3238 2430 3290
rect 2430 3238 2442 3290
rect 2442 3238 2472 3290
rect 2496 3238 2506 3290
rect 2506 3238 2552 3290
rect 2256 3236 2312 3238
rect 2336 3236 2392 3238
rect 2416 3236 2472 3238
rect 2496 3236 2552 3238
rect 4256 4378 4312 4380
rect 4336 4378 4392 4380
rect 4416 4378 4472 4380
rect 4496 4378 4552 4380
rect 4256 4326 4302 4378
rect 4302 4326 4312 4378
rect 4336 4326 4366 4378
rect 4366 4326 4378 4378
rect 4378 4326 4392 4378
rect 4416 4326 4430 4378
rect 4430 4326 4442 4378
rect 4442 4326 4472 4378
rect 4496 4326 4506 4378
rect 4506 4326 4552 4378
rect 4256 4324 4312 4326
rect 4336 4324 4392 4326
rect 4416 4324 4472 4326
rect 4496 4324 4552 4326
rect 3556 3834 3612 3836
rect 3636 3834 3692 3836
rect 3716 3834 3772 3836
rect 3796 3834 3852 3836
rect 3556 3782 3602 3834
rect 3602 3782 3612 3834
rect 3636 3782 3666 3834
rect 3666 3782 3678 3834
rect 3678 3782 3692 3834
rect 3716 3782 3730 3834
rect 3730 3782 3742 3834
rect 3742 3782 3772 3834
rect 3796 3782 3806 3834
rect 3806 3782 3852 3834
rect 3556 3780 3612 3782
rect 3636 3780 3692 3782
rect 3716 3780 3772 3782
rect 3796 3780 3852 3782
rect 1556 2746 1612 2748
rect 1636 2746 1692 2748
rect 1716 2746 1772 2748
rect 1796 2746 1852 2748
rect 1556 2694 1602 2746
rect 1602 2694 1612 2746
rect 1636 2694 1666 2746
rect 1666 2694 1678 2746
rect 1678 2694 1692 2746
rect 1716 2694 1730 2746
rect 1730 2694 1742 2746
rect 1742 2694 1772 2746
rect 1796 2694 1806 2746
rect 1806 2694 1852 2746
rect 1556 2692 1612 2694
rect 1636 2692 1692 2694
rect 1716 2692 1772 2694
rect 1796 2692 1852 2694
rect 3556 2746 3612 2748
rect 3636 2746 3692 2748
rect 3716 2746 3772 2748
rect 3796 2746 3852 2748
rect 3556 2694 3602 2746
rect 3602 2694 3612 2746
rect 3636 2694 3666 2746
rect 3666 2694 3678 2746
rect 3678 2694 3692 2746
rect 3716 2694 3730 2746
rect 3730 2694 3742 2746
rect 3742 2694 3772 2746
rect 3796 2694 3806 2746
rect 3806 2694 3852 2746
rect 3556 2692 3612 2694
rect 3636 2692 3692 2694
rect 3716 2692 3772 2694
rect 3796 2692 3852 2694
rect 4256 3290 4312 3292
rect 4336 3290 4392 3292
rect 4416 3290 4472 3292
rect 4496 3290 4552 3292
rect 4256 3238 4302 3290
rect 4302 3238 4312 3290
rect 4336 3238 4366 3290
rect 4366 3238 4378 3290
rect 4378 3238 4392 3290
rect 4416 3238 4430 3290
rect 4430 3238 4442 3290
rect 4442 3238 4472 3290
rect 4496 3238 4506 3290
rect 4506 3238 4552 3290
rect 4256 3236 4312 3238
rect 4336 3236 4392 3238
rect 4416 3236 4472 3238
rect 4496 3236 4552 3238
rect 5556 6010 5612 6012
rect 5636 6010 5692 6012
rect 5716 6010 5772 6012
rect 5796 6010 5852 6012
rect 5556 5958 5602 6010
rect 5602 5958 5612 6010
rect 5636 5958 5666 6010
rect 5666 5958 5678 6010
rect 5678 5958 5692 6010
rect 5716 5958 5730 6010
rect 5730 5958 5742 6010
rect 5742 5958 5772 6010
rect 5796 5958 5806 6010
rect 5806 5958 5852 6010
rect 5556 5956 5612 5958
rect 5636 5956 5692 5958
rect 5716 5956 5772 5958
rect 5796 5956 5852 5958
rect 6256 5466 6312 5468
rect 6336 5466 6392 5468
rect 6416 5466 6472 5468
rect 6496 5466 6552 5468
rect 6256 5414 6302 5466
rect 6302 5414 6312 5466
rect 6336 5414 6366 5466
rect 6366 5414 6378 5466
rect 6378 5414 6392 5466
rect 6416 5414 6430 5466
rect 6430 5414 6442 5466
rect 6442 5414 6472 5466
rect 6496 5414 6506 5466
rect 6506 5414 6552 5466
rect 6256 5412 6312 5414
rect 6336 5412 6392 5414
rect 6416 5412 6472 5414
rect 6496 5412 6552 5414
rect 5556 4922 5612 4924
rect 5636 4922 5692 4924
rect 5716 4922 5772 4924
rect 5796 4922 5852 4924
rect 5556 4870 5602 4922
rect 5602 4870 5612 4922
rect 5636 4870 5666 4922
rect 5666 4870 5678 4922
rect 5678 4870 5692 4922
rect 5716 4870 5730 4922
rect 5730 4870 5742 4922
rect 5742 4870 5772 4922
rect 5796 4870 5806 4922
rect 5806 4870 5852 4922
rect 5556 4868 5612 4870
rect 5636 4868 5692 4870
rect 5716 4868 5772 4870
rect 5796 4868 5852 4870
rect 5556 3834 5612 3836
rect 5636 3834 5692 3836
rect 5716 3834 5772 3836
rect 5796 3834 5852 3836
rect 5556 3782 5602 3834
rect 5602 3782 5612 3834
rect 5636 3782 5666 3834
rect 5666 3782 5678 3834
rect 5678 3782 5692 3834
rect 5716 3782 5730 3834
rect 5730 3782 5742 3834
rect 5742 3782 5772 3834
rect 5796 3782 5806 3834
rect 5806 3782 5852 3834
rect 5556 3780 5612 3782
rect 5636 3780 5692 3782
rect 5716 3780 5772 3782
rect 5796 3780 5852 3782
rect 8256 9818 8312 9820
rect 8336 9818 8392 9820
rect 8416 9818 8472 9820
rect 8496 9818 8552 9820
rect 8256 9766 8302 9818
rect 8302 9766 8312 9818
rect 8336 9766 8366 9818
rect 8366 9766 8378 9818
rect 8378 9766 8392 9818
rect 8416 9766 8430 9818
rect 8430 9766 8442 9818
rect 8442 9766 8472 9818
rect 8496 9766 8506 9818
rect 8506 9766 8552 9818
rect 8256 9764 8312 9766
rect 8336 9764 8392 9766
rect 8416 9764 8472 9766
rect 8496 9764 8552 9766
rect 7654 9580 7710 9616
rect 7654 9560 7656 9580
rect 7656 9560 7708 9580
rect 7708 9560 7710 9580
rect 7556 9274 7612 9276
rect 7636 9274 7692 9276
rect 7716 9274 7772 9276
rect 7796 9274 7852 9276
rect 7556 9222 7602 9274
rect 7602 9222 7612 9274
rect 7636 9222 7666 9274
rect 7666 9222 7678 9274
rect 7678 9222 7692 9274
rect 7716 9222 7730 9274
rect 7730 9222 7742 9274
rect 7742 9222 7772 9274
rect 7796 9222 7806 9274
rect 7806 9222 7852 9274
rect 7556 9220 7612 9222
rect 7636 9220 7692 9222
rect 7716 9220 7772 9222
rect 7796 9220 7852 9222
rect 8256 8730 8312 8732
rect 8336 8730 8392 8732
rect 8416 8730 8472 8732
rect 8496 8730 8552 8732
rect 8256 8678 8302 8730
rect 8302 8678 8312 8730
rect 8336 8678 8366 8730
rect 8366 8678 8378 8730
rect 8378 8678 8392 8730
rect 8416 8678 8430 8730
rect 8430 8678 8442 8730
rect 8442 8678 8472 8730
rect 8496 8678 8506 8730
rect 8506 8678 8552 8730
rect 8256 8676 8312 8678
rect 8336 8676 8392 8678
rect 8416 8676 8472 8678
rect 8496 8676 8552 8678
rect 7556 8186 7612 8188
rect 7636 8186 7692 8188
rect 7716 8186 7772 8188
rect 7796 8186 7852 8188
rect 7556 8134 7602 8186
rect 7602 8134 7612 8186
rect 7636 8134 7666 8186
rect 7666 8134 7678 8186
rect 7678 8134 7692 8186
rect 7716 8134 7730 8186
rect 7730 8134 7742 8186
rect 7742 8134 7772 8186
rect 7796 8134 7806 8186
rect 7806 8134 7852 8186
rect 7556 8132 7612 8134
rect 7636 8132 7692 8134
rect 7716 8132 7772 8134
rect 7796 8132 7852 8134
rect 7556 7098 7612 7100
rect 7636 7098 7692 7100
rect 7716 7098 7772 7100
rect 7796 7098 7852 7100
rect 7556 7046 7602 7098
rect 7602 7046 7612 7098
rect 7636 7046 7666 7098
rect 7666 7046 7678 7098
rect 7678 7046 7692 7098
rect 7716 7046 7730 7098
rect 7730 7046 7742 7098
rect 7742 7046 7772 7098
rect 7796 7046 7806 7098
rect 7806 7046 7852 7098
rect 7556 7044 7612 7046
rect 7636 7044 7692 7046
rect 7716 7044 7772 7046
rect 7796 7044 7852 7046
rect 8256 7642 8312 7644
rect 8336 7642 8392 7644
rect 8416 7642 8472 7644
rect 8496 7642 8552 7644
rect 8256 7590 8302 7642
rect 8302 7590 8312 7642
rect 8336 7590 8366 7642
rect 8366 7590 8378 7642
rect 8378 7590 8392 7642
rect 8416 7590 8430 7642
rect 8430 7590 8442 7642
rect 8442 7590 8472 7642
rect 8496 7590 8506 7642
rect 8506 7590 8552 7642
rect 8256 7588 8312 7590
rect 8336 7588 8392 7590
rect 8416 7588 8472 7590
rect 8496 7588 8552 7590
rect 9034 9560 9090 9616
rect 9034 8372 9036 8392
rect 9036 8372 9088 8392
rect 9088 8372 9090 8392
rect 9034 8336 9090 8372
rect 10256 10906 10312 10908
rect 10336 10906 10392 10908
rect 10416 10906 10472 10908
rect 10496 10906 10552 10908
rect 10256 10854 10302 10906
rect 10302 10854 10312 10906
rect 10336 10854 10366 10906
rect 10366 10854 10378 10906
rect 10378 10854 10392 10906
rect 10416 10854 10430 10906
rect 10430 10854 10442 10906
rect 10442 10854 10472 10906
rect 10496 10854 10506 10906
rect 10506 10854 10552 10906
rect 10256 10852 10312 10854
rect 10336 10852 10392 10854
rect 10416 10852 10472 10854
rect 10496 10852 10552 10854
rect 9556 10362 9612 10364
rect 9636 10362 9692 10364
rect 9716 10362 9772 10364
rect 9796 10362 9852 10364
rect 9556 10310 9602 10362
rect 9602 10310 9612 10362
rect 9636 10310 9666 10362
rect 9666 10310 9678 10362
rect 9678 10310 9692 10362
rect 9716 10310 9730 10362
rect 9730 10310 9742 10362
rect 9742 10310 9772 10362
rect 9796 10310 9806 10362
rect 9806 10310 9852 10362
rect 9556 10308 9612 10310
rect 9636 10308 9692 10310
rect 9716 10308 9772 10310
rect 9796 10308 9852 10310
rect 9556 9274 9612 9276
rect 9636 9274 9692 9276
rect 9716 9274 9772 9276
rect 9796 9274 9852 9276
rect 9556 9222 9602 9274
rect 9602 9222 9612 9274
rect 9636 9222 9666 9274
rect 9666 9222 9678 9274
rect 9678 9222 9692 9274
rect 9716 9222 9730 9274
rect 9730 9222 9742 9274
rect 9742 9222 9772 9274
rect 9796 9222 9806 9274
rect 9806 9222 9852 9274
rect 9556 9220 9612 9222
rect 9636 9220 9692 9222
rect 9716 9220 9772 9222
rect 9796 9220 9852 9222
rect 10256 9818 10312 9820
rect 10336 9818 10392 9820
rect 10416 9818 10472 9820
rect 10496 9818 10552 9820
rect 10256 9766 10302 9818
rect 10302 9766 10312 9818
rect 10336 9766 10366 9818
rect 10366 9766 10378 9818
rect 10378 9766 10392 9818
rect 10416 9766 10430 9818
rect 10430 9766 10442 9818
rect 10442 9766 10472 9818
rect 10496 9766 10506 9818
rect 10506 9766 10552 9818
rect 10256 9764 10312 9766
rect 10336 9764 10392 9766
rect 10416 9764 10472 9766
rect 10496 9764 10552 9766
rect 9586 8356 9642 8392
rect 9586 8336 9588 8356
rect 9588 8336 9640 8356
rect 9640 8336 9642 8356
rect 9556 8186 9612 8188
rect 9636 8186 9692 8188
rect 9716 8186 9772 8188
rect 9796 8186 9852 8188
rect 9556 8134 9602 8186
rect 9602 8134 9612 8186
rect 9636 8134 9666 8186
rect 9666 8134 9678 8186
rect 9678 8134 9692 8186
rect 9716 8134 9730 8186
rect 9730 8134 9742 8186
rect 9742 8134 9772 8186
rect 9796 8134 9806 8186
rect 9806 8134 9852 8186
rect 9556 8132 9612 8134
rect 9636 8132 9692 8134
rect 9716 8132 9772 8134
rect 9796 8132 9852 8134
rect 10256 8730 10312 8732
rect 10336 8730 10392 8732
rect 10416 8730 10472 8732
rect 10496 8730 10552 8732
rect 10256 8678 10302 8730
rect 10302 8678 10312 8730
rect 10336 8678 10366 8730
rect 10366 8678 10378 8730
rect 10378 8678 10392 8730
rect 10416 8678 10430 8730
rect 10430 8678 10442 8730
rect 10442 8678 10472 8730
rect 10496 8678 10506 8730
rect 10506 8678 10552 8730
rect 10256 8676 10312 8678
rect 10336 8676 10392 8678
rect 10416 8676 10472 8678
rect 10496 8676 10552 8678
rect 10138 8508 10140 8528
rect 10140 8508 10192 8528
rect 10192 8508 10194 8528
rect 10138 8472 10194 8508
rect 11150 12280 11206 12336
rect 11556 12538 11612 12540
rect 11636 12538 11692 12540
rect 11716 12538 11772 12540
rect 11796 12538 11852 12540
rect 11556 12486 11602 12538
rect 11602 12486 11612 12538
rect 11636 12486 11666 12538
rect 11666 12486 11678 12538
rect 11678 12486 11692 12538
rect 11716 12486 11730 12538
rect 11730 12486 11742 12538
rect 11742 12486 11772 12538
rect 11796 12486 11806 12538
rect 11806 12486 11852 12538
rect 11556 12484 11612 12486
rect 11636 12484 11692 12486
rect 11716 12484 11772 12486
rect 11796 12484 11852 12486
rect 11978 11600 12034 11656
rect 11556 11450 11612 11452
rect 11636 11450 11692 11452
rect 11716 11450 11772 11452
rect 11796 11450 11852 11452
rect 11556 11398 11602 11450
rect 11602 11398 11612 11450
rect 11636 11398 11666 11450
rect 11666 11398 11678 11450
rect 11678 11398 11692 11450
rect 11716 11398 11730 11450
rect 11730 11398 11742 11450
rect 11742 11398 11772 11450
rect 11796 11398 11806 11450
rect 11806 11398 11852 11450
rect 11556 11396 11612 11398
rect 11636 11396 11692 11398
rect 11716 11396 11772 11398
rect 11796 11396 11852 11398
rect 11886 10920 11942 10976
rect 8256 6554 8312 6556
rect 8336 6554 8392 6556
rect 8416 6554 8472 6556
rect 8496 6554 8552 6556
rect 8256 6502 8302 6554
rect 8302 6502 8312 6554
rect 8336 6502 8366 6554
rect 8366 6502 8378 6554
rect 8378 6502 8392 6554
rect 8416 6502 8430 6554
rect 8430 6502 8442 6554
rect 8442 6502 8472 6554
rect 8496 6502 8506 6554
rect 8506 6502 8552 6554
rect 8256 6500 8312 6502
rect 8336 6500 8392 6502
rect 8416 6500 8472 6502
rect 8496 6500 8552 6502
rect 7556 6010 7612 6012
rect 7636 6010 7692 6012
rect 7716 6010 7772 6012
rect 7796 6010 7852 6012
rect 7556 5958 7602 6010
rect 7602 5958 7612 6010
rect 7636 5958 7666 6010
rect 7666 5958 7678 6010
rect 7678 5958 7692 6010
rect 7716 5958 7730 6010
rect 7730 5958 7742 6010
rect 7742 5958 7772 6010
rect 7796 5958 7806 6010
rect 7806 5958 7852 6010
rect 7556 5956 7612 5958
rect 7636 5956 7692 5958
rect 7716 5956 7772 5958
rect 7796 5956 7852 5958
rect 6256 4378 6312 4380
rect 6336 4378 6392 4380
rect 6416 4378 6472 4380
rect 6496 4378 6552 4380
rect 6256 4326 6302 4378
rect 6302 4326 6312 4378
rect 6336 4326 6366 4378
rect 6366 4326 6378 4378
rect 6378 4326 6392 4378
rect 6416 4326 6430 4378
rect 6430 4326 6442 4378
rect 6442 4326 6472 4378
rect 6496 4326 6506 4378
rect 6506 4326 6552 4378
rect 6256 4324 6312 4326
rect 6336 4324 6392 4326
rect 6416 4324 6472 4326
rect 6496 4324 6552 4326
rect 6256 3290 6312 3292
rect 6336 3290 6392 3292
rect 6416 3290 6472 3292
rect 6496 3290 6552 3292
rect 6256 3238 6302 3290
rect 6302 3238 6312 3290
rect 6336 3238 6366 3290
rect 6366 3238 6378 3290
rect 6378 3238 6392 3290
rect 6416 3238 6430 3290
rect 6430 3238 6442 3290
rect 6442 3238 6472 3290
rect 6496 3238 6506 3290
rect 6506 3238 6552 3290
rect 6256 3236 6312 3238
rect 6336 3236 6392 3238
rect 6416 3236 6472 3238
rect 6496 3236 6552 3238
rect 8256 5466 8312 5468
rect 8336 5466 8392 5468
rect 8416 5466 8472 5468
rect 8496 5466 8552 5468
rect 8256 5414 8302 5466
rect 8302 5414 8312 5466
rect 8336 5414 8366 5466
rect 8366 5414 8378 5466
rect 8378 5414 8392 5466
rect 8416 5414 8430 5466
rect 8430 5414 8442 5466
rect 8442 5414 8472 5466
rect 8496 5414 8506 5466
rect 8506 5414 8552 5466
rect 8256 5412 8312 5414
rect 8336 5412 8392 5414
rect 8416 5412 8472 5414
rect 8496 5412 8552 5414
rect 7556 4922 7612 4924
rect 7636 4922 7692 4924
rect 7716 4922 7772 4924
rect 7796 4922 7852 4924
rect 7556 4870 7602 4922
rect 7602 4870 7612 4922
rect 7636 4870 7666 4922
rect 7666 4870 7678 4922
rect 7678 4870 7692 4922
rect 7716 4870 7730 4922
rect 7730 4870 7742 4922
rect 7742 4870 7772 4922
rect 7796 4870 7806 4922
rect 7806 4870 7852 4922
rect 7556 4868 7612 4870
rect 7636 4868 7692 4870
rect 7716 4868 7772 4870
rect 7796 4868 7852 4870
rect 5556 2746 5612 2748
rect 5636 2746 5692 2748
rect 5716 2746 5772 2748
rect 5796 2746 5852 2748
rect 5556 2694 5602 2746
rect 5602 2694 5612 2746
rect 5636 2694 5666 2746
rect 5666 2694 5678 2746
rect 5678 2694 5692 2746
rect 5716 2694 5730 2746
rect 5730 2694 5742 2746
rect 5742 2694 5772 2746
rect 5796 2694 5806 2746
rect 5806 2694 5852 2746
rect 5556 2692 5612 2694
rect 5636 2692 5692 2694
rect 5716 2692 5772 2694
rect 5796 2692 5852 2694
rect 7556 3834 7612 3836
rect 7636 3834 7692 3836
rect 7716 3834 7772 3836
rect 7796 3834 7852 3836
rect 7556 3782 7602 3834
rect 7602 3782 7612 3834
rect 7636 3782 7666 3834
rect 7666 3782 7678 3834
rect 7678 3782 7692 3834
rect 7716 3782 7730 3834
rect 7730 3782 7742 3834
rect 7742 3782 7772 3834
rect 7796 3782 7806 3834
rect 7806 3782 7852 3834
rect 7556 3780 7612 3782
rect 7636 3780 7692 3782
rect 7716 3780 7772 3782
rect 7796 3780 7852 3782
rect 8256 4378 8312 4380
rect 8336 4378 8392 4380
rect 8416 4378 8472 4380
rect 8496 4378 8552 4380
rect 8256 4326 8302 4378
rect 8302 4326 8312 4378
rect 8336 4326 8366 4378
rect 8366 4326 8378 4378
rect 8378 4326 8392 4378
rect 8416 4326 8430 4378
rect 8430 4326 8442 4378
rect 8442 4326 8472 4378
rect 8496 4326 8506 4378
rect 8506 4326 8552 4378
rect 8256 4324 8312 4326
rect 8336 4324 8392 4326
rect 8416 4324 8472 4326
rect 8496 4324 8552 4326
rect 9556 7098 9612 7100
rect 9636 7098 9692 7100
rect 9716 7098 9772 7100
rect 9796 7098 9852 7100
rect 9556 7046 9602 7098
rect 9602 7046 9612 7098
rect 9636 7046 9666 7098
rect 9666 7046 9678 7098
rect 9678 7046 9692 7098
rect 9716 7046 9730 7098
rect 9730 7046 9742 7098
rect 9742 7046 9772 7098
rect 9796 7046 9806 7098
rect 9806 7046 9852 7098
rect 9556 7044 9612 7046
rect 9636 7044 9692 7046
rect 9716 7044 9772 7046
rect 9796 7044 9852 7046
rect 11556 10362 11612 10364
rect 11636 10362 11692 10364
rect 11716 10362 11772 10364
rect 11796 10362 11852 10364
rect 11556 10310 11602 10362
rect 11602 10310 11612 10362
rect 11636 10310 11666 10362
rect 11666 10310 11678 10362
rect 11678 10310 11692 10362
rect 11716 10310 11730 10362
rect 11730 10310 11742 10362
rect 11742 10310 11772 10362
rect 11796 10310 11806 10362
rect 11806 10310 11852 10362
rect 11556 10308 11612 10310
rect 11636 10308 11692 10310
rect 11716 10308 11772 10310
rect 11796 10308 11852 10310
rect 11978 10260 12034 10296
rect 11978 10240 11980 10260
rect 11980 10240 12032 10260
rect 12032 10240 12034 10260
rect 11334 8472 11390 8528
rect 12070 9560 12126 9616
rect 11556 9274 11612 9276
rect 11636 9274 11692 9276
rect 11716 9274 11772 9276
rect 11796 9274 11852 9276
rect 11556 9222 11602 9274
rect 11602 9222 11612 9274
rect 11636 9222 11666 9274
rect 11666 9222 11678 9274
rect 11678 9222 11692 9274
rect 11716 9222 11730 9274
rect 11730 9222 11742 9274
rect 11742 9222 11772 9274
rect 11796 9222 11806 9274
rect 11806 9222 11852 9274
rect 11556 9220 11612 9222
rect 11636 9220 11692 9222
rect 11716 9220 11772 9222
rect 11796 9220 11852 9222
rect 11886 8880 11942 8936
rect 11556 8186 11612 8188
rect 11636 8186 11692 8188
rect 11716 8186 11772 8188
rect 11796 8186 11852 8188
rect 11556 8134 11602 8186
rect 11602 8134 11612 8186
rect 11636 8134 11666 8186
rect 11666 8134 11678 8186
rect 11678 8134 11692 8186
rect 11716 8134 11730 8186
rect 11730 8134 11742 8186
rect 11742 8134 11772 8186
rect 11796 8134 11806 8186
rect 11806 8134 11852 8186
rect 11556 8132 11612 8134
rect 11636 8132 11692 8134
rect 11716 8132 11772 8134
rect 11796 8132 11852 8134
rect 12070 8200 12126 8256
rect 10256 7642 10312 7644
rect 10336 7642 10392 7644
rect 10416 7642 10472 7644
rect 10496 7642 10552 7644
rect 10256 7590 10302 7642
rect 10302 7590 10312 7642
rect 10336 7590 10366 7642
rect 10366 7590 10378 7642
rect 10378 7590 10392 7642
rect 10416 7590 10430 7642
rect 10430 7590 10442 7642
rect 10442 7590 10472 7642
rect 10496 7590 10506 7642
rect 10506 7590 10552 7642
rect 10256 7588 10312 7590
rect 10336 7588 10392 7590
rect 10416 7588 10472 7590
rect 10496 7588 10552 7590
rect 9556 6010 9612 6012
rect 9636 6010 9692 6012
rect 9716 6010 9772 6012
rect 9796 6010 9852 6012
rect 9556 5958 9602 6010
rect 9602 5958 9612 6010
rect 9636 5958 9666 6010
rect 9666 5958 9678 6010
rect 9678 5958 9692 6010
rect 9716 5958 9730 6010
rect 9730 5958 9742 6010
rect 9742 5958 9772 6010
rect 9796 5958 9806 6010
rect 9806 5958 9852 6010
rect 9556 5956 9612 5958
rect 9636 5956 9692 5958
rect 9716 5956 9772 5958
rect 9796 5956 9852 5958
rect 9556 4922 9612 4924
rect 9636 4922 9692 4924
rect 9716 4922 9772 4924
rect 9796 4922 9852 4924
rect 9556 4870 9602 4922
rect 9602 4870 9612 4922
rect 9636 4870 9666 4922
rect 9666 4870 9678 4922
rect 9678 4870 9692 4922
rect 9716 4870 9730 4922
rect 9730 4870 9742 4922
rect 9742 4870 9772 4922
rect 9796 4870 9806 4922
rect 9806 4870 9852 4922
rect 9556 4868 9612 4870
rect 9636 4868 9692 4870
rect 9716 4868 9772 4870
rect 9796 4868 9852 4870
rect 10256 6554 10312 6556
rect 10336 6554 10392 6556
rect 10416 6554 10472 6556
rect 10496 6554 10552 6556
rect 10256 6502 10302 6554
rect 10302 6502 10312 6554
rect 10336 6502 10366 6554
rect 10366 6502 10378 6554
rect 10378 6502 10392 6554
rect 10416 6502 10430 6554
rect 10430 6502 10442 6554
rect 10442 6502 10472 6554
rect 10496 6502 10506 6554
rect 10506 6502 10552 6554
rect 10256 6500 10312 6502
rect 10336 6500 10392 6502
rect 10416 6500 10472 6502
rect 10496 6500 10552 6502
rect 10256 5466 10312 5468
rect 10336 5466 10392 5468
rect 10416 5466 10472 5468
rect 10496 5466 10552 5468
rect 10256 5414 10302 5466
rect 10302 5414 10312 5466
rect 10336 5414 10366 5466
rect 10366 5414 10378 5466
rect 10378 5414 10392 5466
rect 10416 5414 10430 5466
rect 10430 5414 10442 5466
rect 10442 5414 10472 5466
rect 10496 5414 10506 5466
rect 10506 5414 10552 5466
rect 10256 5412 10312 5414
rect 10336 5412 10392 5414
rect 10416 5412 10472 5414
rect 10496 5412 10552 5414
rect 7556 2746 7612 2748
rect 7636 2746 7692 2748
rect 7716 2746 7772 2748
rect 7796 2746 7852 2748
rect 7556 2694 7602 2746
rect 7602 2694 7612 2746
rect 7636 2694 7666 2746
rect 7666 2694 7678 2746
rect 7678 2694 7692 2746
rect 7716 2694 7730 2746
rect 7730 2694 7742 2746
rect 7742 2694 7772 2746
rect 7796 2694 7806 2746
rect 7806 2694 7852 2746
rect 7556 2692 7612 2694
rect 7636 2692 7692 2694
rect 7716 2692 7772 2694
rect 7796 2692 7852 2694
rect 8256 3290 8312 3292
rect 8336 3290 8392 3292
rect 8416 3290 8472 3292
rect 8496 3290 8552 3292
rect 8256 3238 8302 3290
rect 8302 3238 8312 3290
rect 8336 3238 8366 3290
rect 8366 3238 8378 3290
rect 8378 3238 8392 3290
rect 8416 3238 8430 3290
rect 8430 3238 8442 3290
rect 8442 3238 8472 3290
rect 8496 3238 8506 3290
rect 8506 3238 8552 3290
rect 8256 3236 8312 3238
rect 8336 3236 8392 3238
rect 8416 3236 8472 3238
rect 8496 3236 8552 3238
rect 9556 3834 9612 3836
rect 9636 3834 9692 3836
rect 9716 3834 9772 3836
rect 9796 3834 9852 3836
rect 9556 3782 9602 3834
rect 9602 3782 9612 3834
rect 9636 3782 9666 3834
rect 9666 3782 9678 3834
rect 9678 3782 9692 3834
rect 9716 3782 9730 3834
rect 9730 3782 9742 3834
rect 9742 3782 9772 3834
rect 9796 3782 9806 3834
rect 9806 3782 9852 3834
rect 9556 3780 9612 3782
rect 9636 3780 9692 3782
rect 9716 3780 9772 3782
rect 9796 3780 9852 3782
rect 11426 7520 11482 7576
rect 11556 7098 11612 7100
rect 11636 7098 11692 7100
rect 11716 7098 11772 7100
rect 11796 7098 11852 7100
rect 11556 7046 11602 7098
rect 11602 7046 11612 7098
rect 11636 7046 11666 7098
rect 11666 7046 11678 7098
rect 11678 7046 11692 7098
rect 11716 7046 11730 7098
rect 11730 7046 11742 7098
rect 11742 7046 11772 7098
rect 11796 7046 11806 7098
rect 11806 7046 11852 7098
rect 11556 7044 11612 7046
rect 11636 7044 11692 7046
rect 11716 7044 11772 7046
rect 11796 7044 11852 7046
rect 11886 6840 11942 6896
rect 10256 4378 10312 4380
rect 10336 4378 10392 4380
rect 10416 4378 10472 4380
rect 10496 4378 10552 4380
rect 10256 4326 10302 4378
rect 10302 4326 10312 4378
rect 10336 4326 10366 4378
rect 10366 4326 10378 4378
rect 10378 4326 10392 4378
rect 10416 4326 10430 4378
rect 10430 4326 10442 4378
rect 10442 4326 10472 4378
rect 10496 4326 10506 4378
rect 10506 4326 10552 4378
rect 10256 4324 10312 4326
rect 10336 4324 10392 4326
rect 10416 4324 10472 4326
rect 10496 4324 10552 4326
rect 10256 3290 10312 3292
rect 10336 3290 10392 3292
rect 10416 3290 10472 3292
rect 10496 3290 10552 3292
rect 10256 3238 10302 3290
rect 10302 3238 10312 3290
rect 10336 3238 10366 3290
rect 10366 3238 10378 3290
rect 10378 3238 10392 3290
rect 10416 3238 10430 3290
rect 10430 3238 10442 3290
rect 10442 3238 10472 3290
rect 10496 3238 10506 3290
rect 10506 3238 10552 3290
rect 10256 3236 10312 3238
rect 10336 3236 10392 3238
rect 10416 3236 10472 3238
rect 10496 3236 10552 3238
rect 9556 2746 9612 2748
rect 9636 2746 9692 2748
rect 9716 2746 9772 2748
rect 9796 2746 9852 2748
rect 9556 2694 9602 2746
rect 9602 2694 9612 2746
rect 9636 2694 9666 2746
rect 9666 2694 9678 2746
rect 9678 2694 9692 2746
rect 9716 2694 9730 2746
rect 9730 2694 9742 2746
rect 9742 2694 9772 2746
rect 9796 2694 9806 2746
rect 9806 2694 9852 2746
rect 9556 2692 9612 2694
rect 9636 2692 9692 2694
rect 9716 2692 9772 2694
rect 9796 2692 9852 2694
rect 11886 6160 11942 6216
rect 11556 6010 11612 6012
rect 11636 6010 11692 6012
rect 11716 6010 11772 6012
rect 11796 6010 11852 6012
rect 11556 5958 11602 6010
rect 11602 5958 11612 6010
rect 11636 5958 11666 6010
rect 11666 5958 11678 6010
rect 11678 5958 11692 6010
rect 11716 5958 11730 6010
rect 11730 5958 11742 6010
rect 11742 5958 11772 6010
rect 11796 5958 11806 6010
rect 11806 5958 11852 6010
rect 11556 5956 11612 5958
rect 11636 5956 11692 5958
rect 11716 5956 11772 5958
rect 11796 5956 11852 5958
rect 11556 4922 11612 4924
rect 11636 4922 11692 4924
rect 11716 4922 11772 4924
rect 11796 4922 11852 4924
rect 11556 4870 11602 4922
rect 11602 4870 11612 4922
rect 11636 4870 11666 4922
rect 11666 4870 11678 4922
rect 11678 4870 11692 4922
rect 11716 4870 11730 4922
rect 11730 4870 11742 4922
rect 11742 4870 11772 4922
rect 11796 4870 11806 4922
rect 11806 4870 11852 4922
rect 11556 4868 11612 4870
rect 11636 4868 11692 4870
rect 11716 4868 11772 4870
rect 11796 4868 11852 4870
rect 12070 5480 12126 5536
rect 11978 4800 12034 4856
rect 11794 4120 11850 4176
rect 11556 3834 11612 3836
rect 11636 3834 11692 3836
rect 11716 3834 11772 3836
rect 11796 3834 11852 3836
rect 11556 3782 11602 3834
rect 11602 3782 11612 3834
rect 11636 3782 11666 3834
rect 11666 3782 11678 3834
rect 11678 3782 11692 3834
rect 11716 3782 11730 3834
rect 11730 3782 11742 3834
rect 11742 3782 11772 3834
rect 11796 3782 11806 3834
rect 11806 3782 11852 3834
rect 11556 3780 11612 3782
rect 11636 3780 11692 3782
rect 11716 3780 11772 3782
rect 11796 3780 11852 3782
rect 11794 3440 11850 3496
rect 11978 2760 12034 2816
rect 11556 2746 11612 2748
rect 11636 2746 11692 2748
rect 11716 2746 11772 2748
rect 11796 2746 11852 2748
rect 11556 2694 11602 2746
rect 11602 2694 11612 2746
rect 11636 2694 11666 2746
rect 11666 2694 11678 2746
rect 11678 2694 11692 2746
rect 11716 2694 11730 2746
rect 11730 2694 11742 2746
rect 11742 2694 11772 2746
rect 11796 2694 11806 2746
rect 11806 2694 11852 2746
rect 11556 2692 11612 2694
rect 11636 2692 11692 2694
rect 11716 2692 11772 2694
rect 11796 2692 11852 2694
rect 2256 2202 2312 2204
rect 2336 2202 2392 2204
rect 2416 2202 2472 2204
rect 2496 2202 2552 2204
rect 2256 2150 2302 2202
rect 2302 2150 2312 2202
rect 2336 2150 2366 2202
rect 2366 2150 2378 2202
rect 2378 2150 2392 2202
rect 2416 2150 2430 2202
rect 2430 2150 2442 2202
rect 2442 2150 2472 2202
rect 2496 2150 2506 2202
rect 2506 2150 2552 2202
rect 2256 2148 2312 2150
rect 2336 2148 2392 2150
rect 2416 2148 2472 2150
rect 2496 2148 2552 2150
rect 4256 2202 4312 2204
rect 4336 2202 4392 2204
rect 4416 2202 4472 2204
rect 4496 2202 4552 2204
rect 4256 2150 4302 2202
rect 4302 2150 4312 2202
rect 4336 2150 4366 2202
rect 4366 2150 4378 2202
rect 4378 2150 4392 2202
rect 4416 2150 4430 2202
rect 4430 2150 4442 2202
rect 4442 2150 4472 2202
rect 4496 2150 4506 2202
rect 4506 2150 4552 2202
rect 4256 2148 4312 2150
rect 4336 2148 4392 2150
rect 4416 2148 4472 2150
rect 4496 2148 4552 2150
rect 6256 2202 6312 2204
rect 6336 2202 6392 2204
rect 6416 2202 6472 2204
rect 6496 2202 6552 2204
rect 6256 2150 6302 2202
rect 6302 2150 6312 2202
rect 6336 2150 6366 2202
rect 6366 2150 6378 2202
rect 6378 2150 6392 2202
rect 6416 2150 6430 2202
rect 6430 2150 6442 2202
rect 6442 2150 6472 2202
rect 6496 2150 6506 2202
rect 6506 2150 6552 2202
rect 6256 2148 6312 2150
rect 6336 2148 6392 2150
rect 6416 2148 6472 2150
rect 6496 2148 6552 2150
rect 8256 2202 8312 2204
rect 8336 2202 8392 2204
rect 8416 2202 8472 2204
rect 8496 2202 8552 2204
rect 8256 2150 8302 2202
rect 8302 2150 8312 2202
rect 8336 2150 8366 2202
rect 8366 2150 8378 2202
rect 8378 2150 8392 2202
rect 8416 2150 8430 2202
rect 8430 2150 8442 2202
rect 8442 2150 8472 2202
rect 8496 2150 8506 2202
rect 8506 2150 8552 2202
rect 8256 2148 8312 2150
rect 8336 2148 8392 2150
rect 8416 2148 8472 2150
rect 8496 2148 8552 2150
rect 10256 2202 10312 2204
rect 10336 2202 10392 2204
rect 10416 2202 10472 2204
rect 10496 2202 10552 2204
rect 10256 2150 10302 2202
rect 10302 2150 10312 2202
rect 10336 2150 10366 2202
rect 10366 2150 10378 2202
rect 10378 2150 10392 2202
rect 10416 2150 10430 2202
rect 10430 2150 10442 2202
rect 10442 2150 10472 2202
rect 10496 2150 10506 2202
rect 10506 2150 10552 2202
rect 10256 2148 10312 2150
rect 10336 2148 10392 2150
rect 10416 2148 10472 2150
rect 10496 2148 10552 2150
<< metal3 >>
rect 2246 13088 2562 13089
rect 2246 13024 2252 13088
rect 2316 13024 2332 13088
rect 2396 13024 2412 13088
rect 2476 13024 2492 13088
rect 2556 13024 2562 13088
rect 2246 13023 2562 13024
rect 4246 13088 4562 13089
rect 4246 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4562 13088
rect 4246 13023 4562 13024
rect 6246 13088 6562 13089
rect 6246 13024 6252 13088
rect 6316 13024 6332 13088
rect 6396 13024 6412 13088
rect 6476 13024 6492 13088
rect 6556 13024 6562 13088
rect 6246 13023 6562 13024
rect 8246 13088 8562 13089
rect 8246 13024 8252 13088
rect 8316 13024 8332 13088
rect 8396 13024 8412 13088
rect 8476 13024 8492 13088
rect 8556 13024 8562 13088
rect 8246 13023 8562 13024
rect 10246 13088 10562 13089
rect 10246 13024 10252 13088
rect 10316 13024 10332 13088
rect 10396 13024 10412 13088
rect 10476 13024 10492 13088
rect 10556 13024 10562 13088
rect 10246 13023 10562 13024
rect 10777 13018 10843 13021
rect 12607 13018 13407 13048
rect 10777 13016 13407 13018
rect 10777 12960 10782 13016
rect 10838 12960 13407 13016
rect 10777 12958 13407 12960
rect 10777 12955 10843 12958
rect 12607 12928 13407 12958
rect 1546 12544 1862 12545
rect 1546 12480 1552 12544
rect 1616 12480 1632 12544
rect 1696 12480 1712 12544
rect 1776 12480 1792 12544
rect 1856 12480 1862 12544
rect 1546 12479 1862 12480
rect 3546 12544 3862 12545
rect 3546 12480 3552 12544
rect 3616 12480 3632 12544
rect 3696 12480 3712 12544
rect 3776 12480 3792 12544
rect 3856 12480 3862 12544
rect 3546 12479 3862 12480
rect 5546 12544 5862 12545
rect 5546 12480 5552 12544
rect 5616 12480 5632 12544
rect 5696 12480 5712 12544
rect 5776 12480 5792 12544
rect 5856 12480 5862 12544
rect 5546 12479 5862 12480
rect 7546 12544 7862 12545
rect 7546 12480 7552 12544
rect 7616 12480 7632 12544
rect 7696 12480 7712 12544
rect 7776 12480 7792 12544
rect 7856 12480 7862 12544
rect 7546 12479 7862 12480
rect 9546 12544 9862 12545
rect 9546 12480 9552 12544
rect 9616 12480 9632 12544
rect 9696 12480 9712 12544
rect 9776 12480 9792 12544
rect 9856 12480 9862 12544
rect 9546 12479 9862 12480
rect 11546 12544 11862 12545
rect 11546 12480 11552 12544
rect 11616 12480 11632 12544
rect 11696 12480 11712 12544
rect 11776 12480 11792 12544
rect 11856 12480 11862 12544
rect 11546 12479 11862 12480
rect 11145 12338 11211 12341
rect 12607 12338 13407 12368
rect 11145 12336 13407 12338
rect 11145 12280 11150 12336
rect 11206 12280 13407 12336
rect 11145 12278 13407 12280
rect 11145 12275 11211 12278
rect 12607 12248 13407 12278
rect 2246 12000 2562 12001
rect 2246 11936 2252 12000
rect 2316 11936 2332 12000
rect 2396 11936 2412 12000
rect 2476 11936 2492 12000
rect 2556 11936 2562 12000
rect 2246 11935 2562 11936
rect 4246 12000 4562 12001
rect 4246 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4562 12000
rect 4246 11935 4562 11936
rect 6246 12000 6562 12001
rect 6246 11936 6252 12000
rect 6316 11936 6332 12000
rect 6396 11936 6412 12000
rect 6476 11936 6492 12000
rect 6556 11936 6562 12000
rect 6246 11935 6562 11936
rect 8246 12000 8562 12001
rect 8246 11936 8252 12000
rect 8316 11936 8332 12000
rect 8396 11936 8412 12000
rect 8476 11936 8492 12000
rect 8556 11936 8562 12000
rect 8246 11935 8562 11936
rect 10246 12000 10562 12001
rect 10246 11936 10252 12000
rect 10316 11936 10332 12000
rect 10396 11936 10412 12000
rect 10476 11936 10492 12000
rect 10556 11936 10562 12000
rect 10246 11935 10562 11936
rect 0 11658 800 11688
rect 4153 11658 4219 11661
rect 0 11656 4219 11658
rect 0 11600 4158 11656
rect 4214 11600 4219 11656
rect 0 11598 4219 11600
rect 0 11568 800 11598
rect 4153 11595 4219 11598
rect 11973 11658 12039 11661
rect 12607 11658 13407 11688
rect 11973 11656 13407 11658
rect 11973 11600 11978 11656
rect 12034 11600 13407 11656
rect 11973 11598 13407 11600
rect 11973 11595 12039 11598
rect 12607 11568 13407 11598
rect 1546 11456 1862 11457
rect 1546 11392 1552 11456
rect 1616 11392 1632 11456
rect 1696 11392 1712 11456
rect 1776 11392 1792 11456
rect 1856 11392 1862 11456
rect 1546 11391 1862 11392
rect 3546 11456 3862 11457
rect 3546 11392 3552 11456
rect 3616 11392 3632 11456
rect 3696 11392 3712 11456
rect 3776 11392 3792 11456
rect 3856 11392 3862 11456
rect 3546 11391 3862 11392
rect 5546 11456 5862 11457
rect 5546 11392 5552 11456
rect 5616 11392 5632 11456
rect 5696 11392 5712 11456
rect 5776 11392 5792 11456
rect 5856 11392 5862 11456
rect 5546 11391 5862 11392
rect 7546 11456 7862 11457
rect 7546 11392 7552 11456
rect 7616 11392 7632 11456
rect 7696 11392 7712 11456
rect 7776 11392 7792 11456
rect 7856 11392 7862 11456
rect 7546 11391 7862 11392
rect 9546 11456 9862 11457
rect 9546 11392 9552 11456
rect 9616 11392 9632 11456
rect 9696 11392 9712 11456
rect 9776 11392 9792 11456
rect 9856 11392 9862 11456
rect 9546 11391 9862 11392
rect 11546 11456 11862 11457
rect 11546 11392 11552 11456
rect 11616 11392 11632 11456
rect 11696 11392 11712 11456
rect 11776 11392 11792 11456
rect 11856 11392 11862 11456
rect 11546 11391 11862 11392
rect 11881 10978 11947 10981
rect 12607 10978 13407 11008
rect 11881 10976 13407 10978
rect 11881 10920 11886 10976
rect 11942 10920 13407 10976
rect 11881 10918 13407 10920
rect 11881 10915 11947 10918
rect 2246 10912 2562 10913
rect 2246 10848 2252 10912
rect 2316 10848 2332 10912
rect 2396 10848 2412 10912
rect 2476 10848 2492 10912
rect 2556 10848 2562 10912
rect 2246 10847 2562 10848
rect 4246 10912 4562 10913
rect 4246 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4562 10912
rect 4246 10847 4562 10848
rect 6246 10912 6562 10913
rect 6246 10848 6252 10912
rect 6316 10848 6332 10912
rect 6396 10848 6412 10912
rect 6476 10848 6492 10912
rect 6556 10848 6562 10912
rect 6246 10847 6562 10848
rect 8246 10912 8562 10913
rect 8246 10848 8252 10912
rect 8316 10848 8332 10912
rect 8396 10848 8412 10912
rect 8476 10848 8492 10912
rect 8556 10848 8562 10912
rect 8246 10847 8562 10848
rect 10246 10912 10562 10913
rect 10246 10848 10252 10912
rect 10316 10848 10332 10912
rect 10396 10848 10412 10912
rect 10476 10848 10492 10912
rect 10556 10848 10562 10912
rect 12607 10888 13407 10918
rect 10246 10847 10562 10848
rect 1546 10368 1862 10369
rect 1546 10304 1552 10368
rect 1616 10304 1632 10368
rect 1696 10304 1712 10368
rect 1776 10304 1792 10368
rect 1856 10304 1862 10368
rect 1546 10303 1862 10304
rect 3546 10368 3862 10369
rect 3546 10304 3552 10368
rect 3616 10304 3632 10368
rect 3696 10304 3712 10368
rect 3776 10304 3792 10368
rect 3856 10304 3862 10368
rect 3546 10303 3862 10304
rect 5546 10368 5862 10369
rect 5546 10304 5552 10368
rect 5616 10304 5632 10368
rect 5696 10304 5712 10368
rect 5776 10304 5792 10368
rect 5856 10304 5862 10368
rect 5546 10303 5862 10304
rect 7546 10368 7862 10369
rect 7546 10304 7552 10368
rect 7616 10304 7632 10368
rect 7696 10304 7712 10368
rect 7776 10304 7792 10368
rect 7856 10304 7862 10368
rect 7546 10303 7862 10304
rect 9546 10368 9862 10369
rect 9546 10304 9552 10368
rect 9616 10304 9632 10368
rect 9696 10304 9712 10368
rect 9776 10304 9792 10368
rect 9856 10304 9862 10368
rect 9546 10303 9862 10304
rect 11546 10368 11862 10369
rect 11546 10304 11552 10368
rect 11616 10304 11632 10368
rect 11696 10304 11712 10368
rect 11776 10304 11792 10368
rect 11856 10304 11862 10368
rect 11546 10303 11862 10304
rect 11973 10298 12039 10301
rect 12607 10298 13407 10328
rect 11973 10296 13407 10298
rect 11973 10240 11978 10296
rect 12034 10240 13407 10296
rect 11973 10238 13407 10240
rect 11973 10235 12039 10238
rect 12607 10208 13407 10238
rect 2246 9824 2562 9825
rect 2246 9760 2252 9824
rect 2316 9760 2332 9824
rect 2396 9760 2412 9824
rect 2476 9760 2492 9824
rect 2556 9760 2562 9824
rect 2246 9759 2562 9760
rect 4246 9824 4562 9825
rect 4246 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4562 9824
rect 4246 9759 4562 9760
rect 6246 9824 6562 9825
rect 6246 9760 6252 9824
rect 6316 9760 6332 9824
rect 6396 9760 6412 9824
rect 6476 9760 6492 9824
rect 6556 9760 6562 9824
rect 6246 9759 6562 9760
rect 8246 9824 8562 9825
rect 8246 9760 8252 9824
rect 8316 9760 8332 9824
rect 8396 9760 8412 9824
rect 8476 9760 8492 9824
rect 8556 9760 8562 9824
rect 8246 9759 8562 9760
rect 10246 9824 10562 9825
rect 10246 9760 10252 9824
rect 10316 9760 10332 9824
rect 10396 9760 10412 9824
rect 10476 9760 10492 9824
rect 10556 9760 10562 9824
rect 10246 9759 10562 9760
rect 0 9618 800 9648
rect 7649 9618 7715 9621
rect 9029 9618 9095 9621
rect 0 9528 858 9618
rect 7649 9616 9095 9618
rect 7649 9560 7654 9616
rect 7710 9560 9034 9616
rect 9090 9560 9095 9616
rect 7649 9558 9095 9560
rect 7649 9555 7715 9558
rect 9029 9555 9095 9558
rect 12065 9618 12131 9621
rect 12607 9618 13407 9648
rect 12065 9616 13407 9618
rect 12065 9560 12070 9616
rect 12126 9560 13407 9616
rect 12065 9558 13407 9560
rect 12065 9555 12131 9558
rect 12607 9528 13407 9558
rect 798 9485 858 9528
rect 798 9480 907 9485
rect 798 9424 846 9480
rect 902 9424 907 9480
rect 798 9422 907 9424
rect 841 9419 907 9422
rect 1546 9280 1862 9281
rect 1546 9216 1552 9280
rect 1616 9216 1632 9280
rect 1696 9216 1712 9280
rect 1776 9216 1792 9280
rect 1856 9216 1862 9280
rect 1546 9215 1862 9216
rect 3546 9280 3862 9281
rect 3546 9216 3552 9280
rect 3616 9216 3632 9280
rect 3696 9216 3712 9280
rect 3776 9216 3792 9280
rect 3856 9216 3862 9280
rect 3546 9215 3862 9216
rect 5546 9280 5862 9281
rect 5546 9216 5552 9280
rect 5616 9216 5632 9280
rect 5696 9216 5712 9280
rect 5776 9216 5792 9280
rect 5856 9216 5862 9280
rect 5546 9215 5862 9216
rect 7546 9280 7862 9281
rect 7546 9216 7552 9280
rect 7616 9216 7632 9280
rect 7696 9216 7712 9280
rect 7776 9216 7792 9280
rect 7856 9216 7862 9280
rect 7546 9215 7862 9216
rect 9546 9280 9862 9281
rect 9546 9216 9552 9280
rect 9616 9216 9632 9280
rect 9696 9216 9712 9280
rect 9776 9216 9792 9280
rect 9856 9216 9862 9280
rect 9546 9215 9862 9216
rect 11546 9280 11862 9281
rect 11546 9216 11552 9280
rect 11616 9216 11632 9280
rect 11696 9216 11712 9280
rect 11776 9216 11792 9280
rect 11856 9216 11862 9280
rect 11546 9215 11862 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 5441 8938 5507 8941
rect 6085 8938 6151 8941
rect 5441 8936 6151 8938
rect 5441 8880 5446 8936
rect 5502 8880 6090 8936
rect 6146 8880 6151 8936
rect 5441 8878 6151 8880
rect 0 8848 800 8878
rect 5441 8875 5507 8878
rect 6085 8875 6151 8878
rect 11881 8938 11947 8941
rect 12607 8938 13407 8968
rect 11881 8936 13407 8938
rect 11881 8880 11886 8936
rect 11942 8880 13407 8936
rect 11881 8878 13407 8880
rect 11881 8875 11947 8878
rect 12607 8848 13407 8878
rect 2246 8736 2562 8737
rect 2246 8672 2252 8736
rect 2316 8672 2332 8736
rect 2396 8672 2412 8736
rect 2476 8672 2492 8736
rect 2556 8672 2562 8736
rect 2246 8671 2562 8672
rect 4246 8736 4562 8737
rect 4246 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4562 8736
rect 4246 8671 4562 8672
rect 6246 8736 6562 8737
rect 6246 8672 6252 8736
rect 6316 8672 6332 8736
rect 6396 8672 6412 8736
rect 6476 8672 6492 8736
rect 6556 8672 6562 8736
rect 6246 8671 6562 8672
rect 8246 8736 8562 8737
rect 8246 8672 8252 8736
rect 8316 8672 8332 8736
rect 8396 8672 8412 8736
rect 8476 8672 8492 8736
rect 8556 8672 8562 8736
rect 8246 8671 8562 8672
rect 10246 8736 10562 8737
rect 10246 8672 10252 8736
rect 10316 8672 10332 8736
rect 10396 8672 10412 8736
rect 10476 8672 10492 8736
rect 10556 8672 10562 8736
rect 10246 8671 10562 8672
rect 10133 8530 10199 8533
rect 11329 8530 11395 8533
rect 10133 8528 11395 8530
rect 10133 8472 10138 8528
rect 10194 8472 11334 8528
rect 11390 8472 11395 8528
rect 10133 8470 11395 8472
rect 10133 8467 10199 8470
rect 11329 8467 11395 8470
rect 9029 8394 9095 8397
rect 9581 8394 9647 8397
rect 9029 8392 9647 8394
rect 9029 8336 9034 8392
rect 9090 8336 9586 8392
rect 9642 8336 9647 8392
rect 9029 8334 9647 8336
rect 9029 8331 9095 8334
rect 9581 8331 9647 8334
rect 0 8258 800 8288
rect 12065 8258 12131 8261
rect 12607 8258 13407 8288
rect 0 8168 858 8258
rect 12065 8256 13407 8258
rect 12065 8200 12070 8256
rect 12126 8200 13407 8256
rect 12065 8198 13407 8200
rect 12065 8195 12131 8198
rect 798 8125 858 8168
rect 1546 8192 1862 8193
rect 1546 8128 1552 8192
rect 1616 8128 1632 8192
rect 1696 8128 1712 8192
rect 1776 8128 1792 8192
rect 1856 8128 1862 8192
rect 1546 8127 1862 8128
rect 3546 8192 3862 8193
rect 3546 8128 3552 8192
rect 3616 8128 3632 8192
rect 3696 8128 3712 8192
rect 3776 8128 3792 8192
rect 3856 8128 3862 8192
rect 3546 8127 3862 8128
rect 5546 8192 5862 8193
rect 5546 8128 5552 8192
rect 5616 8128 5632 8192
rect 5696 8128 5712 8192
rect 5776 8128 5792 8192
rect 5856 8128 5862 8192
rect 5546 8127 5862 8128
rect 7546 8192 7862 8193
rect 7546 8128 7552 8192
rect 7616 8128 7632 8192
rect 7696 8128 7712 8192
rect 7776 8128 7792 8192
rect 7856 8128 7862 8192
rect 7546 8127 7862 8128
rect 9546 8192 9862 8193
rect 9546 8128 9552 8192
rect 9616 8128 9632 8192
rect 9696 8128 9712 8192
rect 9776 8128 9792 8192
rect 9856 8128 9862 8192
rect 9546 8127 9862 8128
rect 11546 8192 11862 8193
rect 11546 8128 11552 8192
rect 11616 8128 11632 8192
rect 11696 8128 11712 8192
rect 11776 8128 11792 8192
rect 11856 8128 11862 8192
rect 12607 8168 13407 8198
rect 11546 8127 11862 8128
rect 798 8120 907 8125
rect 798 8064 846 8120
rect 902 8064 907 8120
rect 798 8062 907 8064
rect 841 8059 907 8062
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 2246 7648 2562 7649
rect 2246 7584 2252 7648
rect 2316 7584 2332 7648
rect 2396 7584 2412 7648
rect 2476 7584 2492 7648
rect 2556 7584 2562 7648
rect 2246 7583 2562 7584
rect 4246 7648 4562 7649
rect 4246 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4562 7648
rect 4246 7583 4562 7584
rect 6246 7648 6562 7649
rect 6246 7584 6252 7648
rect 6316 7584 6332 7648
rect 6396 7584 6412 7648
rect 6476 7584 6492 7648
rect 6556 7584 6562 7648
rect 6246 7583 6562 7584
rect 8246 7648 8562 7649
rect 8246 7584 8252 7648
rect 8316 7584 8332 7648
rect 8396 7584 8412 7648
rect 8476 7584 8492 7648
rect 8556 7584 8562 7648
rect 8246 7583 8562 7584
rect 10246 7648 10562 7649
rect 10246 7584 10252 7648
rect 10316 7584 10332 7648
rect 10396 7584 10412 7648
rect 10476 7584 10492 7648
rect 10556 7584 10562 7648
rect 10246 7583 10562 7584
rect 11421 7578 11487 7581
rect 12607 7578 13407 7608
rect 11421 7576 13407 7578
rect 11421 7520 11426 7576
rect 11482 7520 13407 7576
rect 11421 7518 13407 7520
rect 0 7488 800 7518
rect 11421 7515 11487 7518
rect 12607 7488 13407 7518
rect 1546 7104 1862 7105
rect 1546 7040 1552 7104
rect 1616 7040 1632 7104
rect 1696 7040 1712 7104
rect 1776 7040 1792 7104
rect 1856 7040 1862 7104
rect 1546 7039 1862 7040
rect 3546 7104 3862 7105
rect 3546 7040 3552 7104
rect 3616 7040 3632 7104
rect 3696 7040 3712 7104
rect 3776 7040 3792 7104
rect 3856 7040 3862 7104
rect 3546 7039 3862 7040
rect 5546 7104 5862 7105
rect 5546 7040 5552 7104
rect 5616 7040 5632 7104
rect 5696 7040 5712 7104
rect 5776 7040 5792 7104
rect 5856 7040 5862 7104
rect 5546 7039 5862 7040
rect 7546 7104 7862 7105
rect 7546 7040 7552 7104
rect 7616 7040 7632 7104
rect 7696 7040 7712 7104
rect 7776 7040 7792 7104
rect 7856 7040 7862 7104
rect 7546 7039 7862 7040
rect 9546 7104 9862 7105
rect 9546 7040 9552 7104
rect 9616 7040 9632 7104
rect 9696 7040 9712 7104
rect 9776 7040 9792 7104
rect 9856 7040 9862 7104
rect 9546 7039 9862 7040
rect 11546 7104 11862 7105
rect 11546 7040 11552 7104
rect 11616 7040 11632 7104
rect 11696 7040 11712 7104
rect 11776 7040 11792 7104
rect 11856 7040 11862 7104
rect 11546 7039 11862 7040
rect 11881 6898 11947 6901
rect 12607 6898 13407 6928
rect 11881 6896 13407 6898
rect 11881 6840 11886 6896
rect 11942 6840 13407 6896
rect 11881 6838 13407 6840
rect 11881 6835 11947 6838
rect 12607 6808 13407 6838
rect 2246 6560 2562 6561
rect 2246 6496 2252 6560
rect 2316 6496 2332 6560
rect 2396 6496 2412 6560
rect 2476 6496 2492 6560
rect 2556 6496 2562 6560
rect 2246 6495 2562 6496
rect 4246 6560 4562 6561
rect 4246 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4562 6560
rect 4246 6495 4562 6496
rect 6246 6560 6562 6561
rect 6246 6496 6252 6560
rect 6316 6496 6332 6560
rect 6396 6496 6412 6560
rect 6476 6496 6492 6560
rect 6556 6496 6562 6560
rect 6246 6495 6562 6496
rect 8246 6560 8562 6561
rect 8246 6496 8252 6560
rect 8316 6496 8332 6560
rect 8396 6496 8412 6560
rect 8476 6496 8492 6560
rect 8556 6496 8562 6560
rect 8246 6495 8562 6496
rect 10246 6560 10562 6561
rect 10246 6496 10252 6560
rect 10316 6496 10332 6560
rect 10396 6496 10412 6560
rect 10476 6496 10492 6560
rect 10556 6496 10562 6560
rect 10246 6495 10562 6496
rect 0 6218 800 6248
rect 11881 6218 11947 6221
rect 12607 6218 13407 6248
rect 0 6128 858 6218
rect 11881 6216 13407 6218
rect 11881 6160 11886 6216
rect 11942 6160 13407 6216
rect 11881 6158 13407 6160
rect 11881 6155 11947 6158
rect 12607 6128 13407 6158
rect 798 6085 858 6128
rect 798 6080 907 6085
rect 798 6024 846 6080
rect 902 6024 907 6080
rect 798 6022 907 6024
rect 841 6019 907 6022
rect 1546 6016 1862 6017
rect 1546 5952 1552 6016
rect 1616 5952 1632 6016
rect 1696 5952 1712 6016
rect 1776 5952 1792 6016
rect 1856 5952 1862 6016
rect 1546 5951 1862 5952
rect 3546 6016 3862 6017
rect 3546 5952 3552 6016
rect 3616 5952 3632 6016
rect 3696 5952 3712 6016
rect 3776 5952 3792 6016
rect 3856 5952 3862 6016
rect 3546 5951 3862 5952
rect 5546 6016 5862 6017
rect 5546 5952 5552 6016
rect 5616 5952 5632 6016
rect 5696 5952 5712 6016
rect 5776 5952 5792 6016
rect 5856 5952 5862 6016
rect 5546 5951 5862 5952
rect 7546 6016 7862 6017
rect 7546 5952 7552 6016
rect 7616 5952 7632 6016
rect 7696 5952 7712 6016
rect 7776 5952 7792 6016
rect 7856 5952 7862 6016
rect 7546 5951 7862 5952
rect 9546 6016 9862 6017
rect 9546 5952 9552 6016
rect 9616 5952 9632 6016
rect 9696 5952 9712 6016
rect 9776 5952 9792 6016
rect 9856 5952 9862 6016
rect 9546 5951 9862 5952
rect 11546 6016 11862 6017
rect 11546 5952 11552 6016
rect 11616 5952 11632 6016
rect 11696 5952 11712 6016
rect 11776 5952 11792 6016
rect 11856 5952 11862 6016
rect 11546 5951 11862 5952
rect 0 5538 800 5568
rect 12065 5538 12131 5541
rect 12607 5538 13407 5568
rect 0 5448 858 5538
rect 12065 5536 13407 5538
rect 12065 5480 12070 5536
rect 12126 5480 13407 5536
rect 12065 5478 13407 5480
rect 12065 5475 12131 5478
rect 798 5405 858 5448
rect 2246 5472 2562 5473
rect 2246 5408 2252 5472
rect 2316 5408 2332 5472
rect 2396 5408 2412 5472
rect 2476 5408 2492 5472
rect 2556 5408 2562 5472
rect 2246 5407 2562 5408
rect 4246 5472 4562 5473
rect 4246 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4562 5472
rect 4246 5407 4562 5408
rect 6246 5472 6562 5473
rect 6246 5408 6252 5472
rect 6316 5408 6332 5472
rect 6396 5408 6412 5472
rect 6476 5408 6492 5472
rect 6556 5408 6562 5472
rect 6246 5407 6562 5408
rect 8246 5472 8562 5473
rect 8246 5408 8252 5472
rect 8316 5408 8332 5472
rect 8396 5408 8412 5472
rect 8476 5408 8492 5472
rect 8556 5408 8562 5472
rect 8246 5407 8562 5408
rect 10246 5472 10562 5473
rect 10246 5408 10252 5472
rect 10316 5408 10332 5472
rect 10396 5408 10412 5472
rect 10476 5408 10492 5472
rect 10556 5408 10562 5472
rect 12607 5448 13407 5478
rect 10246 5407 10562 5408
rect 798 5400 907 5405
rect 798 5344 846 5400
rect 902 5344 907 5400
rect 798 5342 907 5344
rect 841 5339 907 5342
rect 1546 4928 1862 4929
rect 1546 4864 1552 4928
rect 1616 4864 1632 4928
rect 1696 4864 1712 4928
rect 1776 4864 1792 4928
rect 1856 4864 1862 4928
rect 1546 4863 1862 4864
rect 3546 4928 3862 4929
rect 3546 4864 3552 4928
rect 3616 4864 3632 4928
rect 3696 4864 3712 4928
rect 3776 4864 3792 4928
rect 3856 4864 3862 4928
rect 3546 4863 3862 4864
rect 5546 4928 5862 4929
rect 5546 4864 5552 4928
rect 5616 4864 5632 4928
rect 5696 4864 5712 4928
rect 5776 4864 5792 4928
rect 5856 4864 5862 4928
rect 5546 4863 5862 4864
rect 7546 4928 7862 4929
rect 7546 4864 7552 4928
rect 7616 4864 7632 4928
rect 7696 4864 7712 4928
rect 7776 4864 7792 4928
rect 7856 4864 7862 4928
rect 7546 4863 7862 4864
rect 9546 4928 9862 4929
rect 9546 4864 9552 4928
rect 9616 4864 9632 4928
rect 9696 4864 9712 4928
rect 9776 4864 9792 4928
rect 9856 4864 9862 4928
rect 9546 4863 9862 4864
rect 11546 4928 11862 4929
rect 11546 4864 11552 4928
rect 11616 4864 11632 4928
rect 11696 4864 11712 4928
rect 11776 4864 11792 4928
rect 11856 4864 11862 4928
rect 11546 4863 11862 4864
rect 11973 4858 12039 4861
rect 12607 4858 13407 4888
rect 11973 4856 13407 4858
rect 11973 4800 11978 4856
rect 12034 4800 13407 4856
rect 11973 4798 13407 4800
rect 11973 4795 12039 4798
rect 12607 4768 13407 4798
rect 2246 4384 2562 4385
rect 2246 4320 2252 4384
rect 2316 4320 2332 4384
rect 2396 4320 2412 4384
rect 2476 4320 2492 4384
rect 2556 4320 2562 4384
rect 2246 4319 2562 4320
rect 4246 4384 4562 4385
rect 4246 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4562 4384
rect 4246 4319 4562 4320
rect 6246 4384 6562 4385
rect 6246 4320 6252 4384
rect 6316 4320 6332 4384
rect 6396 4320 6412 4384
rect 6476 4320 6492 4384
rect 6556 4320 6562 4384
rect 6246 4319 6562 4320
rect 8246 4384 8562 4385
rect 8246 4320 8252 4384
rect 8316 4320 8332 4384
rect 8396 4320 8412 4384
rect 8476 4320 8492 4384
rect 8556 4320 8562 4384
rect 8246 4319 8562 4320
rect 10246 4384 10562 4385
rect 10246 4320 10252 4384
rect 10316 4320 10332 4384
rect 10396 4320 10412 4384
rect 10476 4320 10492 4384
rect 10556 4320 10562 4384
rect 10246 4319 10562 4320
rect 11789 4178 11855 4181
rect 12607 4178 13407 4208
rect 11789 4176 13407 4178
rect 11789 4120 11794 4176
rect 11850 4120 13407 4176
rect 11789 4118 13407 4120
rect 11789 4115 11855 4118
rect 12607 4088 13407 4118
rect 1546 3840 1862 3841
rect 1546 3776 1552 3840
rect 1616 3776 1632 3840
rect 1696 3776 1712 3840
rect 1776 3776 1792 3840
rect 1856 3776 1862 3840
rect 1546 3775 1862 3776
rect 3546 3840 3862 3841
rect 3546 3776 3552 3840
rect 3616 3776 3632 3840
rect 3696 3776 3712 3840
rect 3776 3776 3792 3840
rect 3856 3776 3862 3840
rect 3546 3775 3862 3776
rect 5546 3840 5862 3841
rect 5546 3776 5552 3840
rect 5616 3776 5632 3840
rect 5696 3776 5712 3840
rect 5776 3776 5792 3840
rect 5856 3776 5862 3840
rect 5546 3775 5862 3776
rect 7546 3840 7862 3841
rect 7546 3776 7552 3840
rect 7616 3776 7632 3840
rect 7696 3776 7712 3840
rect 7776 3776 7792 3840
rect 7856 3776 7862 3840
rect 7546 3775 7862 3776
rect 9546 3840 9862 3841
rect 9546 3776 9552 3840
rect 9616 3776 9632 3840
rect 9696 3776 9712 3840
rect 9776 3776 9792 3840
rect 9856 3776 9862 3840
rect 9546 3775 9862 3776
rect 11546 3840 11862 3841
rect 11546 3776 11552 3840
rect 11616 3776 11632 3840
rect 11696 3776 11712 3840
rect 11776 3776 11792 3840
rect 11856 3776 11862 3840
rect 11546 3775 11862 3776
rect 11789 3498 11855 3501
rect 12607 3498 13407 3528
rect 11789 3496 13407 3498
rect 11789 3440 11794 3496
rect 11850 3440 13407 3496
rect 11789 3438 13407 3440
rect 11789 3435 11855 3438
rect 12607 3408 13407 3438
rect 2246 3296 2562 3297
rect 2246 3232 2252 3296
rect 2316 3232 2332 3296
rect 2396 3232 2412 3296
rect 2476 3232 2492 3296
rect 2556 3232 2562 3296
rect 2246 3231 2562 3232
rect 4246 3296 4562 3297
rect 4246 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4562 3296
rect 4246 3231 4562 3232
rect 6246 3296 6562 3297
rect 6246 3232 6252 3296
rect 6316 3232 6332 3296
rect 6396 3232 6412 3296
rect 6476 3232 6492 3296
rect 6556 3232 6562 3296
rect 6246 3231 6562 3232
rect 8246 3296 8562 3297
rect 8246 3232 8252 3296
rect 8316 3232 8332 3296
rect 8396 3232 8412 3296
rect 8476 3232 8492 3296
rect 8556 3232 8562 3296
rect 8246 3231 8562 3232
rect 10246 3296 10562 3297
rect 10246 3232 10252 3296
rect 10316 3232 10332 3296
rect 10396 3232 10412 3296
rect 10476 3232 10492 3296
rect 10556 3232 10562 3296
rect 10246 3231 10562 3232
rect 11973 2818 12039 2821
rect 12607 2818 13407 2848
rect 11973 2816 13407 2818
rect 11973 2760 11978 2816
rect 12034 2760 13407 2816
rect 11973 2758 13407 2760
rect 11973 2755 12039 2758
rect 1546 2752 1862 2753
rect 1546 2688 1552 2752
rect 1616 2688 1632 2752
rect 1696 2688 1712 2752
rect 1776 2688 1792 2752
rect 1856 2688 1862 2752
rect 1546 2687 1862 2688
rect 3546 2752 3862 2753
rect 3546 2688 3552 2752
rect 3616 2688 3632 2752
rect 3696 2688 3712 2752
rect 3776 2688 3792 2752
rect 3856 2688 3862 2752
rect 3546 2687 3862 2688
rect 5546 2752 5862 2753
rect 5546 2688 5552 2752
rect 5616 2688 5632 2752
rect 5696 2688 5712 2752
rect 5776 2688 5792 2752
rect 5856 2688 5862 2752
rect 5546 2687 5862 2688
rect 7546 2752 7862 2753
rect 7546 2688 7552 2752
rect 7616 2688 7632 2752
rect 7696 2688 7712 2752
rect 7776 2688 7792 2752
rect 7856 2688 7862 2752
rect 7546 2687 7862 2688
rect 9546 2752 9862 2753
rect 9546 2688 9552 2752
rect 9616 2688 9632 2752
rect 9696 2688 9712 2752
rect 9776 2688 9792 2752
rect 9856 2688 9862 2752
rect 9546 2687 9862 2688
rect 11546 2752 11862 2753
rect 11546 2688 11552 2752
rect 11616 2688 11632 2752
rect 11696 2688 11712 2752
rect 11776 2688 11792 2752
rect 11856 2688 11862 2752
rect 12607 2728 13407 2758
rect 11546 2687 11862 2688
rect 2246 2208 2562 2209
rect 2246 2144 2252 2208
rect 2316 2144 2332 2208
rect 2396 2144 2412 2208
rect 2476 2144 2492 2208
rect 2556 2144 2562 2208
rect 2246 2143 2562 2144
rect 4246 2208 4562 2209
rect 4246 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4562 2208
rect 4246 2143 4562 2144
rect 6246 2208 6562 2209
rect 6246 2144 6252 2208
rect 6316 2144 6332 2208
rect 6396 2144 6412 2208
rect 6476 2144 6492 2208
rect 6556 2144 6562 2208
rect 6246 2143 6562 2144
rect 8246 2208 8562 2209
rect 8246 2144 8252 2208
rect 8316 2144 8332 2208
rect 8396 2144 8412 2208
rect 8476 2144 8492 2208
rect 8556 2144 8562 2208
rect 8246 2143 8562 2144
rect 10246 2208 10562 2209
rect 10246 2144 10252 2208
rect 10316 2144 10332 2208
rect 10396 2144 10412 2208
rect 10476 2144 10492 2208
rect 10556 2144 10562 2208
rect 10246 2143 10562 2144
<< via3 >>
rect 2252 13084 2316 13088
rect 2252 13028 2256 13084
rect 2256 13028 2312 13084
rect 2312 13028 2316 13084
rect 2252 13024 2316 13028
rect 2332 13084 2396 13088
rect 2332 13028 2336 13084
rect 2336 13028 2392 13084
rect 2392 13028 2396 13084
rect 2332 13024 2396 13028
rect 2412 13084 2476 13088
rect 2412 13028 2416 13084
rect 2416 13028 2472 13084
rect 2472 13028 2476 13084
rect 2412 13024 2476 13028
rect 2492 13084 2556 13088
rect 2492 13028 2496 13084
rect 2496 13028 2552 13084
rect 2552 13028 2556 13084
rect 2492 13024 2556 13028
rect 4252 13084 4316 13088
rect 4252 13028 4256 13084
rect 4256 13028 4312 13084
rect 4312 13028 4316 13084
rect 4252 13024 4316 13028
rect 4332 13084 4396 13088
rect 4332 13028 4336 13084
rect 4336 13028 4392 13084
rect 4392 13028 4396 13084
rect 4332 13024 4396 13028
rect 4412 13084 4476 13088
rect 4412 13028 4416 13084
rect 4416 13028 4472 13084
rect 4472 13028 4476 13084
rect 4412 13024 4476 13028
rect 4492 13084 4556 13088
rect 4492 13028 4496 13084
rect 4496 13028 4552 13084
rect 4552 13028 4556 13084
rect 4492 13024 4556 13028
rect 6252 13084 6316 13088
rect 6252 13028 6256 13084
rect 6256 13028 6312 13084
rect 6312 13028 6316 13084
rect 6252 13024 6316 13028
rect 6332 13084 6396 13088
rect 6332 13028 6336 13084
rect 6336 13028 6392 13084
rect 6392 13028 6396 13084
rect 6332 13024 6396 13028
rect 6412 13084 6476 13088
rect 6412 13028 6416 13084
rect 6416 13028 6472 13084
rect 6472 13028 6476 13084
rect 6412 13024 6476 13028
rect 6492 13084 6556 13088
rect 6492 13028 6496 13084
rect 6496 13028 6552 13084
rect 6552 13028 6556 13084
rect 6492 13024 6556 13028
rect 8252 13084 8316 13088
rect 8252 13028 8256 13084
rect 8256 13028 8312 13084
rect 8312 13028 8316 13084
rect 8252 13024 8316 13028
rect 8332 13084 8396 13088
rect 8332 13028 8336 13084
rect 8336 13028 8392 13084
rect 8392 13028 8396 13084
rect 8332 13024 8396 13028
rect 8412 13084 8476 13088
rect 8412 13028 8416 13084
rect 8416 13028 8472 13084
rect 8472 13028 8476 13084
rect 8412 13024 8476 13028
rect 8492 13084 8556 13088
rect 8492 13028 8496 13084
rect 8496 13028 8552 13084
rect 8552 13028 8556 13084
rect 8492 13024 8556 13028
rect 10252 13084 10316 13088
rect 10252 13028 10256 13084
rect 10256 13028 10312 13084
rect 10312 13028 10316 13084
rect 10252 13024 10316 13028
rect 10332 13084 10396 13088
rect 10332 13028 10336 13084
rect 10336 13028 10392 13084
rect 10392 13028 10396 13084
rect 10332 13024 10396 13028
rect 10412 13084 10476 13088
rect 10412 13028 10416 13084
rect 10416 13028 10472 13084
rect 10472 13028 10476 13084
rect 10412 13024 10476 13028
rect 10492 13084 10556 13088
rect 10492 13028 10496 13084
rect 10496 13028 10552 13084
rect 10552 13028 10556 13084
rect 10492 13024 10556 13028
rect 1552 12540 1616 12544
rect 1552 12484 1556 12540
rect 1556 12484 1612 12540
rect 1612 12484 1616 12540
rect 1552 12480 1616 12484
rect 1632 12540 1696 12544
rect 1632 12484 1636 12540
rect 1636 12484 1692 12540
rect 1692 12484 1696 12540
rect 1632 12480 1696 12484
rect 1712 12540 1776 12544
rect 1712 12484 1716 12540
rect 1716 12484 1772 12540
rect 1772 12484 1776 12540
rect 1712 12480 1776 12484
rect 1792 12540 1856 12544
rect 1792 12484 1796 12540
rect 1796 12484 1852 12540
rect 1852 12484 1856 12540
rect 1792 12480 1856 12484
rect 3552 12540 3616 12544
rect 3552 12484 3556 12540
rect 3556 12484 3612 12540
rect 3612 12484 3616 12540
rect 3552 12480 3616 12484
rect 3632 12540 3696 12544
rect 3632 12484 3636 12540
rect 3636 12484 3692 12540
rect 3692 12484 3696 12540
rect 3632 12480 3696 12484
rect 3712 12540 3776 12544
rect 3712 12484 3716 12540
rect 3716 12484 3772 12540
rect 3772 12484 3776 12540
rect 3712 12480 3776 12484
rect 3792 12540 3856 12544
rect 3792 12484 3796 12540
rect 3796 12484 3852 12540
rect 3852 12484 3856 12540
rect 3792 12480 3856 12484
rect 5552 12540 5616 12544
rect 5552 12484 5556 12540
rect 5556 12484 5612 12540
rect 5612 12484 5616 12540
rect 5552 12480 5616 12484
rect 5632 12540 5696 12544
rect 5632 12484 5636 12540
rect 5636 12484 5692 12540
rect 5692 12484 5696 12540
rect 5632 12480 5696 12484
rect 5712 12540 5776 12544
rect 5712 12484 5716 12540
rect 5716 12484 5772 12540
rect 5772 12484 5776 12540
rect 5712 12480 5776 12484
rect 5792 12540 5856 12544
rect 5792 12484 5796 12540
rect 5796 12484 5852 12540
rect 5852 12484 5856 12540
rect 5792 12480 5856 12484
rect 7552 12540 7616 12544
rect 7552 12484 7556 12540
rect 7556 12484 7612 12540
rect 7612 12484 7616 12540
rect 7552 12480 7616 12484
rect 7632 12540 7696 12544
rect 7632 12484 7636 12540
rect 7636 12484 7692 12540
rect 7692 12484 7696 12540
rect 7632 12480 7696 12484
rect 7712 12540 7776 12544
rect 7712 12484 7716 12540
rect 7716 12484 7772 12540
rect 7772 12484 7776 12540
rect 7712 12480 7776 12484
rect 7792 12540 7856 12544
rect 7792 12484 7796 12540
rect 7796 12484 7852 12540
rect 7852 12484 7856 12540
rect 7792 12480 7856 12484
rect 9552 12540 9616 12544
rect 9552 12484 9556 12540
rect 9556 12484 9612 12540
rect 9612 12484 9616 12540
rect 9552 12480 9616 12484
rect 9632 12540 9696 12544
rect 9632 12484 9636 12540
rect 9636 12484 9692 12540
rect 9692 12484 9696 12540
rect 9632 12480 9696 12484
rect 9712 12540 9776 12544
rect 9712 12484 9716 12540
rect 9716 12484 9772 12540
rect 9772 12484 9776 12540
rect 9712 12480 9776 12484
rect 9792 12540 9856 12544
rect 9792 12484 9796 12540
rect 9796 12484 9852 12540
rect 9852 12484 9856 12540
rect 9792 12480 9856 12484
rect 11552 12540 11616 12544
rect 11552 12484 11556 12540
rect 11556 12484 11612 12540
rect 11612 12484 11616 12540
rect 11552 12480 11616 12484
rect 11632 12540 11696 12544
rect 11632 12484 11636 12540
rect 11636 12484 11692 12540
rect 11692 12484 11696 12540
rect 11632 12480 11696 12484
rect 11712 12540 11776 12544
rect 11712 12484 11716 12540
rect 11716 12484 11772 12540
rect 11772 12484 11776 12540
rect 11712 12480 11776 12484
rect 11792 12540 11856 12544
rect 11792 12484 11796 12540
rect 11796 12484 11852 12540
rect 11852 12484 11856 12540
rect 11792 12480 11856 12484
rect 2252 11996 2316 12000
rect 2252 11940 2256 11996
rect 2256 11940 2312 11996
rect 2312 11940 2316 11996
rect 2252 11936 2316 11940
rect 2332 11996 2396 12000
rect 2332 11940 2336 11996
rect 2336 11940 2392 11996
rect 2392 11940 2396 11996
rect 2332 11936 2396 11940
rect 2412 11996 2476 12000
rect 2412 11940 2416 11996
rect 2416 11940 2472 11996
rect 2472 11940 2476 11996
rect 2412 11936 2476 11940
rect 2492 11996 2556 12000
rect 2492 11940 2496 11996
rect 2496 11940 2552 11996
rect 2552 11940 2556 11996
rect 2492 11936 2556 11940
rect 4252 11996 4316 12000
rect 4252 11940 4256 11996
rect 4256 11940 4312 11996
rect 4312 11940 4316 11996
rect 4252 11936 4316 11940
rect 4332 11996 4396 12000
rect 4332 11940 4336 11996
rect 4336 11940 4392 11996
rect 4392 11940 4396 11996
rect 4332 11936 4396 11940
rect 4412 11996 4476 12000
rect 4412 11940 4416 11996
rect 4416 11940 4472 11996
rect 4472 11940 4476 11996
rect 4412 11936 4476 11940
rect 4492 11996 4556 12000
rect 4492 11940 4496 11996
rect 4496 11940 4552 11996
rect 4552 11940 4556 11996
rect 4492 11936 4556 11940
rect 6252 11996 6316 12000
rect 6252 11940 6256 11996
rect 6256 11940 6312 11996
rect 6312 11940 6316 11996
rect 6252 11936 6316 11940
rect 6332 11996 6396 12000
rect 6332 11940 6336 11996
rect 6336 11940 6392 11996
rect 6392 11940 6396 11996
rect 6332 11936 6396 11940
rect 6412 11996 6476 12000
rect 6412 11940 6416 11996
rect 6416 11940 6472 11996
rect 6472 11940 6476 11996
rect 6412 11936 6476 11940
rect 6492 11996 6556 12000
rect 6492 11940 6496 11996
rect 6496 11940 6552 11996
rect 6552 11940 6556 11996
rect 6492 11936 6556 11940
rect 8252 11996 8316 12000
rect 8252 11940 8256 11996
rect 8256 11940 8312 11996
rect 8312 11940 8316 11996
rect 8252 11936 8316 11940
rect 8332 11996 8396 12000
rect 8332 11940 8336 11996
rect 8336 11940 8392 11996
rect 8392 11940 8396 11996
rect 8332 11936 8396 11940
rect 8412 11996 8476 12000
rect 8412 11940 8416 11996
rect 8416 11940 8472 11996
rect 8472 11940 8476 11996
rect 8412 11936 8476 11940
rect 8492 11996 8556 12000
rect 8492 11940 8496 11996
rect 8496 11940 8552 11996
rect 8552 11940 8556 11996
rect 8492 11936 8556 11940
rect 10252 11996 10316 12000
rect 10252 11940 10256 11996
rect 10256 11940 10312 11996
rect 10312 11940 10316 11996
rect 10252 11936 10316 11940
rect 10332 11996 10396 12000
rect 10332 11940 10336 11996
rect 10336 11940 10392 11996
rect 10392 11940 10396 11996
rect 10332 11936 10396 11940
rect 10412 11996 10476 12000
rect 10412 11940 10416 11996
rect 10416 11940 10472 11996
rect 10472 11940 10476 11996
rect 10412 11936 10476 11940
rect 10492 11996 10556 12000
rect 10492 11940 10496 11996
rect 10496 11940 10552 11996
rect 10552 11940 10556 11996
rect 10492 11936 10556 11940
rect 1552 11452 1616 11456
rect 1552 11396 1556 11452
rect 1556 11396 1612 11452
rect 1612 11396 1616 11452
rect 1552 11392 1616 11396
rect 1632 11452 1696 11456
rect 1632 11396 1636 11452
rect 1636 11396 1692 11452
rect 1692 11396 1696 11452
rect 1632 11392 1696 11396
rect 1712 11452 1776 11456
rect 1712 11396 1716 11452
rect 1716 11396 1772 11452
rect 1772 11396 1776 11452
rect 1712 11392 1776 11396
rect 1792 11452 1856 11456
rect 1792 11396 1796 11452
rect 1796 11396 1852 11452
rect 1852 11396 1856 11452
rect 1792 11392 1856 11396
rect 3552 11452 3616 11456
rect 3552 11396 3556 11452
rect 3556 11396 3612 11452
rect 3612 11396 3616 11452
rect 3552 11392 3616 11396
rect 3632 11452 3696 11456
rect 3632 11396 3636 11452
rect 3636 11396 3692 11452
rect 3692 11396 3696 11452
rect 3632 11392 3696 11396
rect 3712 11452 3776 11456
rect 3712 11396 3716 11452
rect 3716 11396 3772 11452
rect 3772 11396 3776 11452
rect 3712 11392 3776 11396
rect 3792 11452 3856 11456
rect 3792 11396 3796 11452
rect 3796 11396 3852 11452
rect 3852 11396 3856 11452
rect 3792 11392 3856 11396
rect 5552 11452 5616 11456
rect 5552 11396 5556 11452
rect 5556 11396 5612 11452
rect 5612 11396 5616 11452
rect 5552 11392 5616 11396
rect 5632 11452 5696 11456
rect 5632 11396 5636 11452
rect 5636 11396 5692 11452
rect 5692 11396 5696 11452
rect 5632 11392 5696 11396
rect 5712 11452 5776 11456
rect 5712 11396 5716 11452
rect 5716 11396 5772 11452
rect 5772 11396 5776 11452
rect 5712 11392 5776 11396
rect 5792 11452 5856 11456
rect 5792 11396 5796 11452
rect 5796 11396 5852 11452
rect 5852 11396 5856 11452
rect 5792 11392 5856 11396
rect 7552 11452 7616 11456
rect 7552 11396 7556 11452
rect 7556 11396 7612 11452
rect 7612 11396 7616 11452
rect 7552 11392 7616 11396
rect 7632 11452 7696 11456
rect 7632 11396 7636 11452
rect 7636 11396 7692 11452
rect 7692 11396 7696 11452
rect 7632 11392 7696 11396
rect 7712 11452 7776 11456
rect 7712 11396 7716 11452
rect 7716 11396 7772 11452
rect 7772 11396 7776 11452
rect 7712 11392 7776 11396
rect 7792 11452 7856 11456
rect 7792 11396 7796 11452
rect 7796 11396 7852 11452
rect 7852 11396 7856 11452
rect 7792 11392 7856 11396
rect 9552 11452 9616 11456
rect 9552 11396 9556 11452
rect 9556 11396 9612 11452
rect 9612 11396 9616 11452
rect 9552 11392 9616 11396
rect 9632 11452 9696 11456
rect 9632 11396 9636 11452
rect 9636 11396 9692 11452
rect 9692 11396 9696 11452
rect 9632 11392 9696 11396
rect 9712 11452 9776 11456
rect 9712 11396 9716 11452
rect 9716 11396 9772 11452
rect 9772 11396 9776 11452
rect 9712 11392 9776 11396
rect 9792 11452 9856 11456
rect 9792 11396 9796 11452
rect 9796 11396 9852 11452
rect 9852 11396 9856 11452
rect 9792 11392 9856 11396
rect 11552 11452 11616 11456
rect 11552 11396 11556 11452
rect 11556 11396 11612 11452
rect 11612 11396 11616 11452
rect 11552 11392 11616 11396
rect 11632 11452 11696 11456
rect 11632 11396 11636 11452
rect 11636 11396 11692 11452
rect 11692 11396 11696 11452
rect 11632 11392 11696 11396
rect 11712 11452 11776 11456
rect 11712 11396 11716 11452
rect 11716 11396 11772 11452
rect 11772 11396 11776 11452
rect 11712 11392 11776 11396
rect 11792 11452 11856 11456
rect 11792 11396 11796 11452
rect 11796 11396 11852 11452
rect 11852 11396 11856 11452
rect 11792 11392 11856 11396
rect 2252 10908 2316 10912
rect 2252 10852 2256 10908
rect 2256 10852 2312 10908
rect 2312 10852 2316 10908
rect 2252 10848 2316 10852
rect 2332 10908 2396 10912
rect 2332 10852 2336 10908
rect 2336 10852 2392 10908
rect 2392 10852 2396 10908
rect 2332 10848 2396 10852
rect 2412 10908 2476 10912
rect 2412 10852 2416 10908
rect 2416 10852 2472 10908
rect 2472 10852 2476 10908
rect 2412 10848 2476 10852
rect 2492 10908 2556 10912
rect 2492 10852 2496 10908
rect 2496 10852 2552 10908
rect 2552 10852 2556 10908
rect 2492 10848 2556 10852
rect 4252 10908 4316 10912
rect 4252 10852 4256 10908
rect 4256 10852 4312 10908
rect 4312 10852 4316 10908
rect 4252 10848 4316 10852
rect 4332 10908 4396 10912
rect 4332 10852 4336 10908
rect 4336 10852 4392 10908
rect 4392 10852 4396 10908
rect 4332 10848 4396 10852
rect 4412 10908 4476 10912
rect 4412 10852 4416 10908
rect 4416 10852 4472 10908
rect 4472 10852 4476 10908
rect 4412 10848 4476 10852
rect 4492 10908 4556 10912
rect 4492 10852 4496 10908
rect 4496 10852 4552 10908
rect 4552 10852 4556 10908
rect 4492 10848 4556 10852
rect 6252 10908 6316 10912
rect 6252 10852 6256 10908
rect 6256 10852 6312 10908
rect 6312 10852 6316 10908
rect 6252 10848 6316 10852
rect 6332 10908 6396 10912
rect 6332 10852 6336 10908
rect 6336 10852 6392 10908
rect 6392 10852 6396 10908
rect 6332 10848 6396 10852
rect 6412 10908 6476 10912
rect 6412 10852 6416 10908
rect 6416 10852 6472 10908
rect 6472 10852 6476 10908
rect 6412 10848 6476 10852
rect 6492 10908 6556 10912
rect 6492 10852 6496 10908
rect 6496 10852 6552 10908
rect 6552 10852 6556 10908
rect 6492 10848 6556 10852
rect 8252 10908 8316 10912
rect 8252 10852 8256 10908
rect 8256 10852 8312 10908
rect 8312 10852 8316 10908
rect 8252 10848 8316 10852
rect 8332 10908 8396 10912
rect 8332 10852 8336 10908
rect 8336 10852 8392 10908
rect 8392 10852 8396 10908
rect 8332 10848 8396 10852
rect 8412 10908 8476 10912
rect 8412 10852 8416 10908
rect 8416 10852 8472 10908
rect 8472 10852 8476 10908
rect 8412 10848 8476 10852
rect 8492 10908 8556 10912
rect 8492 10852 8496 10908
rect 8496 10852 8552 10908
rect 8552 10852 8556 10908
rect 8492 10848 8556 10852
rect 10252 10908 10316 10912
rect 10252 10852 10256 10908
rect 10256 10852 10312 10908
rect 10312 10852 10316 10908
rect 10252 10848 10316 10852
rect 10332 10908 10396 10912
rect 10332 10852 10336 10908
rect 10336 10852 10392 10908
rect 10392 10852 10396 10908
rect 10332 10848 10396 10852
rect 10412 10908 10476 10912
rect 10412 10852 10416 10908
rect 10416 10852 10472 10908
rect 10472 10852 10476 10908
rect 10412 10848 10476 10852
rect 10492 10908 10556 10912
rect 10492 10852 10496 10908
rect 10496 10852 10552 10908
rect 10552 10852 10556 10908
rect 10492 10848 10556 10852
rect 1552 10364 1616 10368
rect 1552 10308 1556 10364
rect 1556 10308 1612 10364
rect 1612 10308 1616 10364
rect 1552 10304 1616 10308
rect 1632 10364 1696 10368
rect 1632 10308 1636 10364
rect 1636 10308 1692 10364
rect 1692 10308 1696 10364
rect 1632 10304 1696 10308
rect 1712 10364 1776 10368
rect 1712 10308 1716 10364
rect 1716 10308 1772 10364
rect 1772 10308 1776 10364
rect 1712 10304 1776 10308
rect 1792 10364 1856 10368
rect 1792 10308 1796 10364
rect 1796 10308 1852 10364
rect 1852 10308 1856 10364
rect 1792 10304 1856 10308
rect 3552 10364 3616 10368
rect 3552 10308 3556 10364
rect 3556 10308 3612 10364
rect 3612 10308 3616 10364
rect 3552 10304 3616 10308
rect 3632 10364 3696 10368
rect 3632 10308 3636 10364
rect 3636 10308 3692 10364
rect 3692 10308 3696 10364
rect 3632 10304 3696 10308
rect 3712 10364 3776 10368
rect 3712 10308 3716 10364
rect 3716 10308 3772 10364
rect 3772 10308 3776 10364
rect 3712 10304 3776 10308
rect 3792 10364 3856 10368
rect 3792 10308 3796 10364
rect 3796 10308 3852 10364
rect 3852 10308 3856 10364
rect 3792 10304 3856 10308
rect 5552 10364 5616 10368
rect 5552 10308 5556 10364
rect 5556 10308 5612 10364
rect 5612 10308 5616 10364
rect 5552 10304 5616 10308
rect 5632 10364 5696 10368
rect 5632 10308 5636 10364
rect 5636 10308 5692 10364
rect 5692 10308 5696 10364
rect 5632 10304 5696 10308
rect 5712 10364 5776 10368
rect 5712 10308 5716 10364
rect 5716 10308 5772 10364
rect 5772 10308 5776 10364
rect 5712 10304 5776 10308
rect 5792 10364 5856 10368
rect 5792 10308 5796 10364
rect 5796 10308 5852 10364
rect 5852 10308 5856 10364
rect 5792 10304 5856 10308
rect 7552 10364 7616 10368
rect 7552 10308 7556 10364
rect 7556 10308 7612 10364
rect 7612 10308 7616 10364
rect 7552 10304 7616 10308
rect 7632 10364 7696 10368
rect 7632 10308 7636 10364
rect 7636 10308 7692 10364
rect 7692 10308 7696 10364
rect 7632 10304 7696 10308
rect 7712 10364 7776 10368
rect 7712 10308 7716 10364
rect 7716 10308 7772 10364
rect 7772 10308 7776 10364
rect 7712 10304 7776 10308
rect 7792 10364 7856 10368
rect 7792 10308 7796 10364
rect 7796 10308 7852 10364
rect 7852 10308 7856 10364
rect 7792 10304 7856 10308
rect 9552 10364 9616 10368
rect 9552 10308 9556 10364
rect 9556 10308 9612 10364
rect 9612 10308 9616 10364
rect 9552 10304 9616 10308
rect 9632 10364 9696 10368
rect 9632 10308 9636 10364
rect 9636 10308 9692 10364
rect 9692 10308 9696 10364
rect 9632 10304 9696 10308
rect 9712 10364 9776 10368
rect 9712 10308 9716 10364
rect 9716 10308 9772 10364
rect 9772 10308 9776 10364
rect 9712 10304 9776 10308
rect 9792 10364 9856 10368
rect 9792 10308 9796 10364
rect 9796 10308 9852 10364
rect 9852 10308 9856 10364
rect 9792 10304 9856 10308
rect 11552 10364 11616 10368
rect 11552 10308 11556 10364
rect 11556 10308 11612 10364
rect 11612 10308 11616 10364
rect 11552 10304 11616 10308
rect 11632 10364 11696 10368
rect 11632 10308 11636 10364
rect 11636 10308 11692 10364
rect 11692 10308 11696 10364
rect 11632 10304 11696 10308
rect 11712 10364 11776 10368
rect 11712 10308 11716 10364
rect 11716 10308 11772 10364
rect 11772 10308 11776 10364
rect 11712 10304 11776 10308
rect 11792 10364 11856 10368
rect 11792 10308 11796 10364
rect 11796 10308 11852 10364
rect 11852 10308 11856 10364
rect 11792 10304 11856 10308
rect 2252 9820 2316 9824
rect 2252 9764 2256 9820
rect 2256 9764 2312 9820
rect 2312 9764 2316 9820
rect 2252 9760 2316 9764
rect 2332 9820 2396 9824
rect 2332 9764 2336 9820
rect 2336 9764 2392 9820
rect 2392 9764 2396 9820
rect 2332 9760 2396 9764
rect 2412 9820 2476 9824
rect 2412 9764 2416 9820
rect 2416 9764 2472 9820
rect 2472 9764 2476 9820
rect 2412 9760 2476 9764
rect 2492 9820 2556 9824
rect 2492 9764 2496 9820
rect 2496 9764 2552 9820
rect 2552 9764 2556 9820
rect 2492 9760 2556 9764
rect 4252 9820 4316 9824
rect 4252 9764 4256 9820
rect 4256 9764 4312 9820
rect 4312 9764 4316 9820
rect 4252 9760 4316 9764
rect 4332 9820 4396 9824
rect 4332 9764 4336 9820
rect 4336 9764 4392 9820
rect 4392 9764 4396 9820
rect 4332 9760 4396 9764
rect 4412 9820 4476 9824
rect 4412 9764 4416 9820
rect 4416 9764 4472 9820
rect 4472 9764 4476 9820
rect 4412 9760 4476 9764
rect 4492 9820 4556 9824
rect 4492 9764 4496 9820
rect 4496 9764 4552 9820
rect 4552 9764 4556 9820
rect 4492 9760 4556 9764
rect 6252 9820 6316 9824
rect 6252 9764 6256 9820
rect 6256 9764 6312 9820
rect 6312 9764 6316 9820
rect 6252 9760 6316 9764
rect 6332 9820 6396 9824
rect 6332 9764 6336 9820
rect 6336 9764 6392 9820
rect 6392 9764 6396 9820
rect 6332 9760 6396 9764
rect 6412 9820 6476 9824
rect 6412 9764 6416 9820
rect 6416 9764 6472 9820
rect 6472 9764 6476 9820
rect 6412 9760 6476 9764
rect 6492 9820 6556 9824
rect 6492 9764 6496 9820
rect 6496 9764 6552 9820
rect 6552 9764 6556 9820
rect 6492 9760 6556 9764
rect 8252 9820 8316 9824
rect 8252 9764 8256 9820
rect 8256 9764 8312 9820
rect 8312 9764 8316 9820
rect 8252 9760 8316 9764
rect 8332 9820 8396 9824
rect 8332 9764 8336 9820
rect 8336 9764 8392 9820
rect 8392 9764 8396 9820
rect 8332 9760 8396 9764
rect 8412 9820 8476 9824
rect 8412 9764 8416 9820
rect 8416 9764 8472 9820
rect 8472 9764 8476 9820
rect 8412 9760 8476 9764
rect 8492 9820 8556 9824
rect 8492 9764 8496 9820
rect 8496 9764 8552 9820
rect 8552 9764 8556 9820
rect 8492 9760 8556 9764
rect 10252 9820 10316 9824
rect 10252 9764 10256 9820
rect 10256 9764 10312 9820
rect 10312 9764 10316 9820
rect 10252 9760 10316 9764
rect 10332 9820 10396 9824
rect 10332 9764 10336 9820
rect 10336 9764 10392 9820
rect 10392 9764 10396 9820
rect 10332 9760 10396 9764
rect 10412 9820 10476 9824
rect 10412 9764 10416 9820
rect 10416 9764 10472 9820
rect 10472 9764 10476 9820
rect 10412 9760 10476 9764
rect 10492 9820 10556 9824
rect 10492 9764 10496 9820
rect 10496 9764 10552 9820
rect 10552 9764 10556 9820
rect 10492 9760 10556 9764
rect 1552 9276 1616 9280
rect 1552 9220 1556 9276
rect 1556 9220 1612 9276
rect 1612 9220 1616 9276
rect 1552 9216 1616 9220
rect 1632 9276 1696 9280
rect 1632 9220 1636 9276
rect 1636 9220 1692 9276
rect 1692 9220 1696 9276
rect 1632 9216 1696 9220
rect 1712 9276 1776 9280
rect 1712 9220 1716 9276
rect 1716 9220 1772 9276
rect 1772 9220 1776 9276
rect 1712 9216 1776 9220
rect 1792 9276 1856 9280
rect 1792 9220 1796 9276
rect 1796 9220 1852 9276
rect 1852 9220 1856 9276
rect 1792 9216 1856 9220
rect 3552 9276 3616 9280
rect 3552 9220 3556 9276
rect 3556 9220 3612 9276
rect 3612 9220 3616 9276
rect 3552 9216 3616 9220
rect 3632 9276 3696 9280
rect 3632 9220 3636 9276
rect 3636 9220 3692 9276
rect 3692 9220 3696 9276
rect 3632 9216 3696 9220
rect 3712 9276 3776 9280
rect 3712 9220 3716 9276
rect 3716 9220 3772 9276
rect 3772 9220 3776 9276
rect 3712 9216 3776 9220
rect 3792 9276 3856 9280
rect 3792 9220 3796 9276
rect 3796 9220 3852 9276
rect 3852 9220 3856 9276
rect 3792 9216 3856 9220
rect 5552 9276 5616 9280
rect 5552 9220 5556 9276
rect 5556 9220 5612 9276
rect 5612 9220 5616 9276
rect 5552 9216 5616 9220
rect 5632 9276 5696 9280
rect 5632 9220 5636 9276
rect 5636 9220 5692 9276
rect 5692 9220 5696 9276
rect 5632 9216 5696 9220
rect 5712 9276 5776 9280
rect 5712 9220 5716 9276
rect 5716 9220 5772 9276
rect 5772 9220 5776 9276
rect 5712 9216 5776 9220
rect 5792 9276 5856 9280
rect 5792 9220 5796 9276
rect 5796 9220 5852 9276
rect 5852 9220 5856 9276
rect 5792 9216 5856 9220
rect 7552 9276 7616 9280
rect 7552 9220 7556 9276
rect 7556 9220 7612 9276
rect 7612 9220 7616 9276
rect 7552 9216 7616 9220
rect 7632 9276 7696 9280
rect 7632 9220 7636 9276
rect 7636 9220 7692 9276
rect 7692 9220 7696 9276
rect 7632 9216 7696 9220
rect 7712 9276 7776 9280
rect 7712 9220 7716 9276
rect 7716 9220 7772 9276
rect 7772 9220 7776 9276
rect 7712 9216 7776 9220
rect 7792 9276 7856 9280
rect 7792 9220 7796 9276
rect 7796 9220 7852 9276
rect 7852 9220 7856 9276
rect 7792 9216 7856 9220
rect 9552 9276 9616 9280
rect 9552 9220 9556 9276
rect 9556 9220 9612 9276
rect 9612 9220 9616 9276
rect 9552 9216 9616 9220
rect 9632 9276 9696 9280
rect 9632 9220 9636 9276
rect 9636 9220 9692 9276
rect 9692 9220 9696 9276
rect 9632 9216 9696 9220
rect 9712 9276 9776 9280
rect 9712 9220 9716 9276
rect 9716 9220 9772 9276
rect 9772 9220 9776 9276
rect 9712 9216 9776 9220
rect 9792 9276 9856 9280
rect 9792 9220 9796 9276
rect 9796 9220 9852 9276
rect 9852 9220 9856 9276
rect 9792 9216 9856 9220
rect 11552 9276 11616 9280
rect 11552 9220 11556 9276
rect 11556 9220 11612 9276
rect 11612 9220 11616 9276
rect 11552 9216 11616 9220
rect 11632 9276 11696 9280
rect 11632 9220 11636 9276
rect 11636 9220 11692 9276
rect 11692 9220 11696 9276
rect 11632 9216 11696 9220
rect 11712 9276 11776 9280
rect 11712 9220 11716 9276
rect 11716 9220 11772 9276
rect 11772 9220 11776 9276
rect 11712 9216 11776 9220
rect 11792 9276 11856 9280
rect 11792 9220 11796 9276
rect 11796 9220 11852 9276
rect 11852 9220 11856 9276
rect 11792 9216 11856 9220
rect 2252 8732 2316 8736
rect 2252 8676 2256 8732
rect 2256 8676 2312 8732
rect 2312 8676 2316 8732
rect 2252 8672 2316 8676
rect 2332 8732 2396 8736
rect 2332 8676 2336 8732
rect 2336 8676 2392 8732
rect 2392 8676 2396 8732
rect 2332 8672 2396 8676
rect 2412 8732 2476 8736
rect 2412 8676 2416 8732
rect 2416 8676 2472 8732
rect 2472 8676 2476 8732
rect 2412 8672 2476 8676
rect 2492 8732 2556 8736
rect 2492 8676 2496 8732
rect 2496 8676 2552 8732
rect 2552 8676 2556 8732
rect 2492 8672 2556 8676
rect 4252 8732 4316 8736
rect 4252 8676 4256 8732
rect 4256 8676 4312 8732
rect 4312 8676 4316 8732
rect 4252 8672 4316 8676
rect 4332 8732 4396 8736
rect 4332 8676 4336 8732
rect 4336 8676 4392 8732
rect 4392 8676 4396 8732
rect 4332 8672 4396 8676
rect 4412 8732 4476 8736
rect 4412 8676 4416 8732
rect 4416 8676 4472 8732
rect 4472 8676 4476 8732
rect 4412 8672 4476 8676
rect 4492 8732 4556 8736
rect 4492 8676 4496 8732
rect 4496 8676 4552 8732
rect 4552 8676 4556 8732
rect 4492 8672 4556 8676
rect 6252 8732 6316 8736
rect 6252 8676 6256 8732
rect 6256 8676 6312 8732
rect 6312 8676 6316 8732
rect 6252 8672 6316 8676
rect 6332 8732 6396 8736
rect 6332 8676 6336 8732
rect 6336 8676 6392 8732
rect 6392 8676 6396 8732
rect 6332 8672 6396 8676
rect 6412 8732 6476 8736
rect 6412 8676 6416 8732
rect 6416 8676 6472 8732
rect 6472 8676 6476 8732
rect 6412 8672 6476 8676
rect 6492 8732 6556 8736
rect 6492 8676 6496 8732
rect 6496 8676 6552 8732
rect 6552 8676 6556 8732
rect 6492 8672 6556 8676
rect 8252 8732 8316 8736
rect 8252 8676 8256 8732
rect 8256 8676 8312 8732
rect 8312 8676 8316 8732
rect 8252 8672 8316 8676
rect 8332 8732 8396 8736
rect 8332 8676 8336 8732
rect 8336 8676 8392 8732
rect 8392 8676 8396 8732
rect 8332 8672 8396 8676
rect 8412 8732 8476 8736
rect 8412 8676 8416 8732
rect 8416 8676 8472 8732
rect 8472 8676 8476 8732
rect 8412 8672 8476 8676
rect 8492 8732 8556 8736
rect 8492 8676 8496 8732
rect 8496 8676 8552 8732
rect 8552 8676 8556 8732
rect 8492 8672 8556 8676
rect 10252 8732 10316 8736
rect 10252 8676 10256 8732
rect 10256 8676 10312 8732
rect 10312 8676 10316 8732
rect 10252 8672 10316 8676
rect 10332 8732 10396 8736
rect 10332 8676 10336 8732
rect 10336 8676 10392 8732
rect 10392 8676 10396 8732
rect 10332 8672 10396 8676
rect 10412 8732 10476 8736
rect 10412 8676 10416 8732
rect 10416 8676 10472 8732
rect 10472 8676 10476 8732
rect 10412 8672 10476 8676
rect 10492 8732 10556 8736
rect 10492 8676 10496 8732
rect 10496 8676 10552 8732
rect 10552 8676 10556 8732
rect 10492 8672 10556 8676
rect 1552 8188 1616 8192
rect 1552 8132 1556 8188
rect 1556 8132 1612 8188
rect 1612 8132 1616 8188
rect 1552 8128 1616 8132
rect 1632 8188 1696 8192
rect 1632 8132 1636 8188
rect 1636 8132 1692 8188
rect 1692 8132 1696 8188
rect 1632 8128 1696 8132
rect 1712 8188 1776 8192
rect 1712 8132 1716 8188
rect 1716 8132 1772 8188
rect 1772 8132 1776 8188
rect 1712 8128 1776 8132
rect 1792 8188 1856 8192
rect 1792 8132 1796 8188
rect 1796 8132 1852 8188
rect 1852 8132 1856 8188
rect 1792 8128 1856 8132
rect 3552 8188 3616 8192
rect 3552 8132 3556 8188
rect 3556 8132 3612 8188
rect 3612 8132 3616 8188
rect 3552 8128 3616 8132
rect 3632 8188 3696 8192
rect 3632 8132 3636 8188
rect 3636 8132 3692 8188
rect 3692 8132 3696 8188
rect 3632 8128 3696 8132
rect 3712 8188 3776 8192
rect 3712 8132 3716 8188
rect 3716 8132 3772 8188
rect 3772 8132 3776 8188
rect 3712 8128 3776 8132
rect 3792 8188 3856 8192
rect 3792 8132 3796 8188
rect 3796 8132 3852 8188
rect 3852 8132 3856 8188
rect 3792 8128 3856 8132
rect 5552 8188 5616 8192
rect 5552 8132 5556 8188
rect 5556 8132 5612 8188
rect 5612 8132 5616 8188
rect 5552 8128 5616 8132
rect 5632 8188 5696 8192
rect 5632 8132 5636 8188
rect 5636 8132 5692 8188
rect 5692 8132 5696 8188
rect 5632 8128 5696 8132
rect 5712 8188 5776 8192
rect 5712 8132 5716 8188
rect 5716 8132 5772 8188
rect 5772 8132 5776 8188
rect 5712 8128 5776 8132
rect 5792 8188 5856 8192
rect 5792 8132 5796 8188
rect 5796 8132 5852 8188
rect 5852 8132 5856 8188
rect 5792 8128 5856 8132
rect 7552 8188 7616 8192
rect 7552 8132 7556 8188
rect 7556 8132 7612 8188
rect 7612 8132 7616 8188
rect 7552 8128 7616 8132
rect 7632 8188 7696 8192
rect 7632 8132 7636 8188
rect 7636 8132 7692 8188
rect 7692 8132 7696 8188
rect 7632 8128 7696 8132
rect 7712 8188 7776 8192
rect 7712 8132 7716 8188
rect 7716 8132 7772 8188
rect 7772 8132 7776 8188
rect 7712 8128 7776 8132
rect 7792 8188 7856 8192
rect 7792 8132 7796 8188
rect 7796 8132 7852 8188
rect 7852 8132 7856 8188
rect 7792 8128 7856 8132
rect 9552 8188 9616 8192
rect 9552 8132 9556 8188
rect 9556 8132 9612 8188
rect 9612 8132 9616 8188
rect 9552 8128 9616 8132
rect 9632 8188 9696 8192
rect 9632 8132 9636 8188
rect 9636 8132 9692 8188
rect 9692 8132 9696 8188
rect 9632 8128 9696 8132
rect 9712 8188 9776 8192
rect 9712 8132 9716 8188
rect 9716 8132 9772 8188
rect 9772 8132 9776 8188
rect 9712 8128 9776 8132
rect 9792 8188 9856 8192
rect 9792 8132 9796 8188
rect 9796 8132 9852 8188
rect 9852 8132 9856 8188
rect 9792 8128 9856 8132
rect 11552 8188 11616 8192
rect 11552 8132 11556 8188
rect 11556 8132 11612 8188
rect 11612 8132 11616 8188
rect 11552 8128 11616 8132
rect 11632 8188 11696 8192
rect 11632 8132 11636 8188
rect 11636 8132 11692 8188
rect 11692 8132 11696 8188
rect 11632 8128 11696 8132
rect 11712 8188 11776 8192
rect 11712 8132 11716 8188
rect 11716 8132 11772 8188
rect 11772 8132 11776 8188
rect 11712 8128 11776 8132
rect 11792 8188 11856 8192
rect 11792 8132 11796 8188
rect 11796 8132 11852 8188
rect 11852 8132 11856 8188
rect 11792 8128 11856 8132
rect 2252 7644 2316 7648
rect 2252 7588 2256 7644
rect 2256 7588 2312 7644
rect 2312 7588 2316 7644
rect 2252 7584 2316 7588
rect 2332 7644 2396 7648
rect 2332 7588 2336 7644
rect 2336 7588 2392 7644
rect 2392 7588 2396 7644
rect 2332 7584 2396 7588
rect 2412 7644 2476 7648
rect 2412 7588 2416 7644
rect 2416 7588 2472 7644
rect 2472 7588 2476 7644
rect 2412 7584 2476 7588
rect 2492 7644 2556 7648
rect 2492 7588 2496 7644
rect 2496 7588 2552 7644
rect 2552 7588 2556 7644
rect 2492 7584 2556 7588
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 4332 7644 4396 7648
rect 4332 7588 4336 7644
rect 4336 7588 4392 7644
rect 4392 7588 4396 7644
rect 4332 7584 4396 7588
rect 4412 7644 4476 7648
rect 4412 7588 4416 7644
rect 4416 7588 4472 7644
rect 4472 7588 4476 7644
rect 4412 7584 4476 7588
rect 4492 7644 4556 7648
rect 4492 7588 4496 7644
rect 4496 7588 4552 7644
rect 4552 7588 4556 7644
rect 4492 7584 4556 7588
rect 6252 7644 6316 7648
rect 6252 7588 6256 7644
rect 6256 7588 6312 7644
rect 6312 7588 6316 7644
rect 6252 7584 6316 7588
rect 6332 7644 6396 7648
rect 6332 7588 6336 7644
rect 6336 7588 6392 7644
rect 6392 7588 6396 7644
rect 6332 7584 6396 7588
rect 6412 7644 6476 7648
rect 6412 7588 6416 7644
rect 6416 7588 6472 7644
rect 6472 7588 6476 7644
rect 6412 7584 6476 7588
rect 6492 7644 6556 7648
rect 6492 7588 6496 7644
rect 6496 7588 6552 7644
rect 6552 7588 6556 7644
rect 6492 7584 6556 7588
rect 8252 7644 8316 7648
rect 8252 7588 8256 7644
rect 8256 7588 8312 7644
rect 8312 7588 8316 7644
rect 8252 7584 8316 7588
rect 8332 7644 8396 7648
rect 8332 7588 8336 7644
rect 8336 7588 8392 7644
rect 8392 7588 8396 7644
rect 8332 7584 8396 7588
rect 8412 7644 8476 7648
rect 8412 7588 8416 7644
rect 8416 7588 8472 7644
rect 8472 7588 8476 7644
rect 8412 7584 8476 7588
rect 8492 7644 8556 7648
rect 8492 7588 8496 7644
rect 8496 7588 8552 7644
rect 8552 7588 8556 7644
rect 8492 7584 8556 7588
rect 10252 7644 10316 7648
rect 10252 7588 10256 7644
rect 10256 7588 10312 7644
rect 10312 7588 10316 7644
rect 10252 7584 10316 7588
rect 10332 7644 10396 7648
rect 10332 7588 10336 7644
rect 10336 7588 10392 7644
rect 10392 7588 10396 7644
rect 10332 7584 10396 7588
rect 10412 7644 10476 7648
rect 10412 7588 10416 7644
rect 10416 7588 10472 7644
rect 10472 7588 10476 7644
rect 10412 7584 10476 7588
rect 10492 7644 10556 7648
rect 10492 7588 10496 7644
rect 10496 7588 10552 7644
rect 10552 7588 10556 7644
rect 10492 7584 10556 7588
rect 1552 7100 1616 7104
rect 1552 7044 1556 7100
rect 1556 7044 1612 7100
rect 1612 7044 1616 7100
rect 1552 7040 1616 7044
rect 1632 7100 1696 7104
rect 1632 7044 1636 7100
rect 1636 7044 1692 7100
rect 1692 7044 1696 7100
rect 1632 7040 1696 7044
rect 1712 7100 1776 7104
rect 1712 7044 1716 7100
rect 1716 7044 1772 7100
rect 1772 7044 1776 7100
rect 1712 7040 1776 7044
rect 1792 7100 1856 7104
rect 1792 7044 1796 7100
rect 1796 7044 1852 7100
rect 1852 7044 1856 7100
rect 1792 7040 1856 7044
rect 3552 7100 3616 7104
rect 3552 7044 3556 7100
rect 3556 7044 3612 7100
rect 3612 7044 3616 7100
rect 3552 7040 3616 7044
rect 3632 7100 3696 7104
rect 3632 7044 3636 7100
rect 3636 7044 3692 7100
rect 3692 7044 3696 7100
rect 3632 7040 3696 7044
rect 3712 7100 3776 7104
rect 3712 7044 3716 7100
rect 3716 7044 3772 7100
rect 3772 7044 3776 7100
rect 3712 7040 3776 7044
rect 3792 7100 3856 7104
rect 3792 7044 3796 7100
rect 3796 7044 3852 7100
rect 3852 7044 3856 7100
rect 3792 7040 3856 7044
rect 5552 7100 5616 7104
rect 5552 7044 5556 7100
rect 5556 7044 5612 7100
rect 5612 7044 5616 7100
rect 5552 7040 5616 7044
rect 5632 7100 5696 7104
rect 5632 7044 5636 7100
rect 5636 7044 5692 7100
rect 5692 7044 5696 7100
rect 5632 7040 5696 7044
rect 5712 7100 5776 7104
rect 5712 7044 5716 7100
rect 5716 7044 5772 7100
rect 5772 7044 5776 7100
rect 5712 7040 5776 7044
rect 5792 7100 5856 7104
rect 5792 7044 5796 7100
rect 5796 7044 5852 7100
rect 5852 7044 5856 7100
rect 5792 7040 5856 7044
rect 7552 7100 7616 7104
rect 7552 7044 7556 7100
rect 7556 7044 7612 7100
rect 7612 7044 7616 7100
rect 7552 7040 7616 7044
rect 7632 7100 7696 7104
rect 7632 7044 7636 7100
rect 7636 7044 7692 7100
rect 7692 7044 7696 7100
rect 7632 7040 7696 7044
rect 7712 7100 7776 7104
rect 7712 7044 7716 7100
rect 7716 7044 7772 7100
rect 7772 7044 7776 7100
rect 7712 7040 7776 7044
rect 7792 7100 7856 7104
rect 7792 7044 7796 7100
rect 7796 7044 7852 7100
rect 7852 7044 7856 7100
rect 7792 7040 7856 7044
rect 9552 7100 9616 7104
rect 9552 7044 9556 7100
rect 9556 7044 9612 7100
rect 9612 7044 9616 7100
rect 9552 7040 9616 7044
rect 9632 7100 9696 7104
rect 9632 7044 9636 7100
rect 9636 7044 9692 7100
rect 9692 7044 9696 7100
rect 9632 7040 9696 7044
rect 9712 7100 9776 7104
rect 9712 7044 9716 7100
rect 9716 7044 9772 7100
rect 9772 7044 9776 7100
rect 9712 7040 9776 7044
rect 9792 7100 9856 7104
rect 9792 7044 9796 7100
rect 9796 7044 9852 7100
rect 9852 7044 9856 7100
rect 9792 7040 9856 7044
rect 11552 7100 11616 7104
rect 11552 7044 11556 7100
rect 11556 7044 11612 7100
rect 11612 7044 11616 7100
rect 11552 7040 11616 7044
rect 11632 7100 11696 7104
rect 11632 7044 11636 7100
rect 11636 7044 11692 7100
rect 11692 7044 11696 7100
rect 11632 7040 11696 7044
rect 11712 7100 11776 7104
rect 11712 7044 11716 7100
rect 11716 7044 11772 7100
rect 11772 7044 11776 7100
rect 11712 7040 11776 7044
rect 11792 7100 11856 7104
rect 11792 7044 11796 7100
rect 11796 7044 11852 7100
rect 11852 7044 11856 7100
rect 11792 7040 11856 7044
rect 2252 6556 2316 6560
rect 2252 6500 2256 6556
rect 2256 6500 2312 6556
rect 2312 6500 2316 6556
rect 2252 6496 2316 6500
rect 2332 6556 2396 6560
rect 2332 6500 2336 6556
rect 2336 6500 2392 6556
rect 2392 6500 2396 6556
rect 2332 6496 2396 6500
rect 2412 6556 2476 6560
rect 2412 6500 2416 6556
rect 2416 6500 2472 6556
rect 2472 6500 2476 6556
rect 2412 6496 2476 6500
rect 2492 6556 2556 6560
rect 2492 6500 2496 6556
rect 2496 6500 2552 6556
rect 2552 6500 2556 6556
rect 2492 6496 2556 6500
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 4332 6556 4396 6560
rect 4332 6500 4336 6556
rect 4336 6500 4392 6556
rect 4392 6500 4396 6556
rect 4332 6496 4396 6500
rect 4412 6556 4476 6560
rect 4412 6500 4416 6556
rect 4416 6500 4472 6556
rect 4472 6500 4476 6556
rect 4412 6496 4476 6500
rect 4492 6556 4556 6560
rect 4492 6500 4496 6556
rect 4496 6500 4552 6556
rect 4552 6500 4556 6556
rect 4492 6496 4556 6500
rect 6252 6556 6316 6560
rect 6252 6500 6256 6556
rect 6256 6500 6312 6556
rect 6312 6500 6316 6556
rect 6252 6496 6316 6500
rect 6332 6556 6396 6560
rect 6332 6500 6336 6556
rect 6336 6500 6392 6556
rect 6392 6500 6396 6556
rect 6332 6496 6396 6500
rect 6412 6556 6476 6560
rect 6412 6500 6416 6556
rect 6416 6500 6472 6556
rect 6472 6500 6476 6556
rect 6412 6496 6476 6500
rect 6492 6556 6556 6560
rect 6492 6500 6496 6556
rect 6496 6500 6552 6556
rect 6552 6500 6556 6556
rect 6492 6496 6556 6500
rect 8252 6556 8316 6560
rect 8252 6500 8256 6556
rect 8256 6500 8312 6556
rect 8312 6500 8316 6556
rect 8252 6496 8316 6500
rect 8332 6556 8396 6560
rect 8332 6500 8336 6556
rect 8336 6500 8392 6556
rect 8392 6500 8396 6556
rect 8332 6496 8396 6500
rect 8412 6556 8476 6560
rect 8412 6500 8416 6556
rect 8416 6500 8472 6556
rect 8472 6500 8476 6556
rect 8412 6496 8476 6500
rect 8492 6556 8556 6560
rect 8492 6500 8496 6556
rect 8496 6500 8552 6556
rect 8552 6500 8556 6556
rect 8492 6496 8556 6500
rect 10252 6556 10316 6560
rect 10252 6500 10256 6556
rect 10256 6500 10312 6556
rect 10312 6500 10316 6556
rect 10252 6496 10316 6500
rect 10332 6556 10396 6560
rect 10332 6500 10336 6556
rect 10336 6500 10392 6556
rect 10392 6500 10396 6556
rect 10332 6496 10396 6500
rect 10412 6556 10476 6560
rect 10412 6500 10416 6556
rect 10416 6500 10472 6556
rect 10472 6500 10476 6556
rect 10412 6496 10476 6500
rect 10492 6556 10556 6560
rect 10492 6500 10496 6556
rect 10496 6500 10552 6556
rect 10552 6500 10556 6556
rect 10492 6496 10556 6500
rect 1552 6012 1616 6016
rect 1552 5956 1556 6012
rect 1556 5956 1612 6012
rect 1612 5956 1616 6012
rect 1552 5952 1616 5956
rect 1632 6012 1696 6016
rect 1632 5956 1636 6012
rect 1636 5956 1692 6012
rect 1692 5956 1696 6012
rect 1632 5952 1696 5956
rect 1712 6012 1776 6016
rect 1712 5956 1716 6012
rect 1716 5956 1772 6012
rect 1772 5956 1776 6012
rect 1712 5952 1776 5956
rect 1792 6012 1856 6016
rect 1792 5956 1796 6012
rect 1796 5956 1852 6012
rect 1852 5956 1856 6012
rect 1792 5952 1856 5956
rect 3552 6012 3616 6016
rect 3552 5956 3556 6012
rect 3556 5956 3612 6012
rect 3612 5956 3616 6012
rect 3552 5952 3616 5956
rect 3632 6012 3696 6016
rect 3632 5956 3636 6012
rect 3636 5956 3692 6012
rect 3692 5956 3696 6012
rect 3632 5952 3696 5956
rect 3712 6012 3776 6016
rect 3712 5956 3716 6012
rect 3716 5956 3772 6012
rect 3772 5956 3776 6012
rect 3712 5952 3776 5956
rect 3792 6012 3856 6016
rect 3792 5956 3796 6012
rect 3796 5956 3852 6012
rect 3852 5956 3856 6012
rect 3792 5952 3856 5956
rect 5552 6012 5616 6016
rect 5552 5956 5556 6012
rect 5556 5956 5612 6012
rect 5612 5956 5616 6012
rect 5552 5952 5616 5956
rect 5632 6012 5696 6016
rect 5632 5956 5636 6012
rect 5636 5956 5692 6012
rect 5692 5956 5696 6012
rect 5632 5952 5696 5956
rect 5712 6012 5776 6016
rect 5712 5956 5716 6012
rect 5716 5956 5772 6012
rect 5772 5956 5776 6012
rect 5712 5952 5776 5956
rect 5792 6012 5856 6016
rect 5792 5956 5796 6012
rect 5796 5956 5852 6012
rect 5852 5956 5856 6012
rect 5792 5952 5856 5956
rect 7552 6012 7616 6016
rect 7552 5956 7556 6012
rect 7556 5956 7612 6012
rect 7612 5956 7616 6012
rect 7552 5952 7616 5956
rect 7632 6012 7696 6016
rect 7632 5956 7636 6012
rect 7636 5956 7692 6012
rect 7692 5956 7696 6012
rect 7632 5952 7696 5956
rect 7712 6012 7776 6016
rect 7712 5956 7716 6012
rect 7716 5956 7772 6012
rect 7772 5956 7776 6012
rect 7712 5952 7776 5956
rect 7792 6012 7856 6016
rect 7792 5956 7796 6012
rect 7796 5956 7852 6012
rect 7852 5956 7856 6012
rect 7792 5952 7856 5956
rect 9552 6012 9616 6016
rect 9552 5956 9556 6012
rect 9556 5956 9612 6012
rect 9612 5956 9616 6012
rect 9552 5952 9616 5956
rect 9632 6012 9696 6016
rect 9632 5956 9636 6012
rect 9636 5956 9692 6012
rect 9692 5956 9696 6012
rect 9632 5952 9696 5956
rect 9712 6012 9776 6016
rect 9712 5956 9716 6012
rect 9716 5956 9772 6012
rect 9772 5956 9776 6012
rect 9712 5952 9776 5956
rect 9792 6012 9856 6016
rect 9792 5956 9796 6012
rect 9796 5956 9852 6012
rect 9852 5956 9856 6012
rect 9792 5952 9856 5956
rect 11552 6012 11616 6016
rect 11552 5956 11556 6012
rect 11556 5956 11612 6012
rect 11612 5956 11616 6012
rect 11552 5952 11616 5956
rect 11632 6012 11696 6016
rect 11632 5956 11636 6012
rect 11636 5956 11692 6012
rect 11692 5956 11696 6012
rect 11632 5952 11696 5956
rect 11712 6012 11776 6016
rect 11712 5956 11716 6012
rect 11716 5956 11772 6012
rect 11772 5956 11776 6012
rect 11712 5952 11776 5956
rect 11792 6012 11856 6016
rect 11792 5956 11796 6012
rect 11796 5956 11852 6012
rect 11852 5956 11856 6012
rect 11792 5952 11856 5956
rect 2252 5468 2316 5472
rect 2252 5412 2256 5468
rect 2256 5412 2312 5468
rect 2312 5412 2316 5468
rect 2252 5408 2316 5412
rect 2332 5468 2396 5472
rect 2332 5412 2336 5468
rect 2336 5412 2392 5468
rect 2392 5412 2396 5468
rect 2332 5408 2396 5412
rect 2412 5468 2476 5472
rect 2412 5412 2416 5468
rect 2416 5412 2472 5468
rect 2472 5412 2476 5468
rect 2412 5408 2476 5412
rect 2492 5468 2556 5472
rect 2492 5412 2496 5468
rect 2496 5412 2552 5468
rect 2552 5412 2556 5468
rect 2492 5408 2556 5412
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 4332 5468 4396 5472
rect 4332 5412 4336 5468
rect 4336 5412 4392 5468
rect 4392 5412 4396 5468
rect 4332 5408 4396 5412
rect 4412 5468 4476 5472
rect 4412 5412 4416 5468
rect 4416 5412 4472 5468
rect 4472 5412 4476 5468
rect 4412 5408 4476 5412
rect 4492 5468 4556 5472
rect 4492 5412 4496 5468
rect 4496 5412 4552 5468
rect 4552 5412 4556 5468
rect 4492 5408 4556 5412
rect 6252 5468 6316 5472
rect 6252 5412 6256 5468
rect 6256 5412 6312 5468
rect 6312 5412 6316 5468
rect 6252 5408 6316 5412
rect 6332 5468 6396 5472
rect 6332 5412 6336 5468
rect 6336 5412 6392 5468
rect 6392 5412 6396 5468
rect 6332 5408 6396 5412
rect 6412 5468 6476 5472
rect 6412 5412 6416 5468
rect 6416 5412 6472 5468
rect 6472 5412 6476 5468
rect 6412 5408 6476 5412
rect 6492 5468 6556 5472
rect 6492 5412 6496 5468
rect 6496 5412 6552 5468
rect 6552 5412 6556 5468
rect 6492 5408 6556 5412
rect 8252 5468 8316 5472
rect 8252 5412 8256 5468
rect 8256 5412 8312 5468
rect 8312 5412 8316 5468
rect 8252 5408 8316 5412
rect 8332 5468 8396 5472
rect 8332 5412 8336 5468
rect 8336 5412 8392 5468
rect 8392 5412 8396 5468
rect 8332 5408 8396 5412
rect 8412 5468 8476 5472
rect 8412 5412 8416 5468
rect 8416 5412 8472 5468
rect 8472 5412 8476 5468
rect 8412 5408 8476 5412
rect 8492 5468 8556 5472
rect 8492 5412 8496 5468
rect 8496 5412 8552 5468
rect 8552 5412 8556 5468
rect 8492 5408 8556 5412
rect 10252 5468 10316 5472
rect 10252 5412 10256 5468
rect 10256 5412 10312 5468
rect 10312 5412 10316 5468
rect 10252 5408 10316 5412
rect 10332 5468 10396 5472
rect 10332 5412 10336 5468
rect 10336 5412 10392 5468
rect 10392 5412 10396 5468
rect 10332 5408 10396 5412
rect 10412 5468 10476 5472
rect 10412 5412 10416 5468
rect 10416 5412 10472 5468
rect 10472 5412 10476 5468
rect 10412 5408 10476 5412
rect 10492 5468 10556 5472
rect 10492 5412 10496 5468
rect 10496 5412 10552 5468
rect 10552 5412 10556 5468
rect 10492 5408 10556 5412
rect 1552 4924 1616 4928
rect 1552 4868 1556 4924
rect 1556 4868 1612 4924
rect 1612 4868 1616 4924
rect 1552 4864 1616 4868
rect 1632 4924 1696 4928
rect 1632 4868 1636 4924
rect 1636 4868 1692 4924
rect 1692 4868 1696 4924
rect 1632 4864 1696 4868
rect 1712 4924 1776 4928
rect 1712 4868 1716 4924
rect 1716 4868 1772 4924
rect 1772 4868 1776 4924
rect 1712 4864 1776 4868
rect 1792 4924 1856 4928
rect 1792 4868 1796 4924
rect 1796 4868 1852 4924
rect 1852 4868 1856 4924
rect 1792 4864 1856 4868
rect 3552 4924 3616 4928
rect 3552 4868 3556 4924
rect 3556 4868 3612 4924
rect 3612 4868 3616 4924
rect 3552 4864 3616 4868
rect 3632 4924 3696 4928
rect 3632 4868 3636 4924
rect 3636 4868 3692 4924
rect 3692 4868 3696 4924
rect 3632 4864 3696 4868
rect 3712 4924 3776 4928
rect 3712 4868 3716 4924
rect 3716 4868 3772 4924
rect 3772 4868 3776 4924
rect 3712 4864 3776 4868
rect 3792 4924 3856 4928
rect 3792 4868 3796 4924
rect 3796 4868 3852 4924
rect 3852 4868 3856 4924
rect 3792 4864 3856 4868
rect 5552 4924 5616 4928
rect 5552 4868 5556 4924
rect 5556 4868 5612 4924
rect 5612 4868 5616 4924
rect 5552 4864 5616 4868
rect 5632 4924 5696 4928
rect 5632 4868 5636 4924
rect 5636 4868 5692 4924
rect 5692 4868 5696 4924
rect 5632 4864 5696 4868
rect 5712 4924 5776 4928
rect 5712 4868 5716 4924
rect 5716 4868 5772 4924
rect 5772 4868 5776 4924
rect 5712 4864 5776 4868
rect 5792 4924 5856 4928
rect 5792 4868 5796 4924
rect 5796 4868 5852 4924
rect 5852 4868 5856 4924
rect 5792 4864 5856 4868
rect 7552 4924 7616 4928
rect 7552 4868 7556 4924
rect 7556 4868 7612 4924
rect 7612 4868 7616 4924
rect 7552 4864 7616 4868
rect 7632 4924 7696 4928
rect 7632 4868 7636 4924
rect 7636 4868 7692 4924
rect 7692 4868 7696 4924
rect 7632 4864 7696 4868
rect 7712 4924 7776 4928
rect 7712 4868 7716 4924
rect 7716 4868 7772 4924
rect 7772 4868 7776 4924
rect 7712 4864 7776 4868
rect 7792 4924 7856 4928
rect 7792 4868 7796 4924
rect 7796 4868 7852 4924
rect 7852 4868 7856 4924
rect 7792 4864 7856 4868
rect 9552 4924 9616 4928
rect 9552 4868 9556 4924
rect 9556 4868 9612 4924
rect 9612 4868 9616 4924
rect 9552 4864 9616 4868
rect 9632 4924 9696 4928
rect 9632 4868 9636 4924
rect 9636 4868 9692 4924
rect 9692 4868 9696 4924
rect 9632 4864 9696 4868
rect 9712 4924 9776 4928
rect 9712 4868 9716 4924
rect 9716 4868 9772 4924
rect 9772 4868 9776 4924
rect 9712 4864 9776 4868
rect 9792 4924 9856 4928
rect 9792 4868 9796 4924
rect 9796 4868 9852 4924
rect 9852 4868 9856 4924
rect 9792 4864 9856 4868
rect 11552 4924 11616 4928
rect 11552 4868 11556 4924
rect 11556 4868 11612 4924
rect 11612 4868 11616 4924
rect 11552 4864 11616 4868
rect 11632 4924 11696 4928
rect 11632 4868 11636 4924
rect 11636 4868 11692 4924
rect 11692 4868 11696 4924
rect 11632 4864 11696 4868
rect 11712 4924 11776 4928
rect 11712 4868 11716 4924
rect 11716 4868 11772 4924
rect 11772 4868 11776 4924
rect 11712 4864 11776 4868
rect 11792 4924 11856 4928
rect 11792 4868 11796 4924
rect 11796 4868 11852 4924
rect 11852 4868 11856 4924
rect 11792 4864 11856 4868
rect 2252 4380 2316 4384
rect 2252 4324 2256 4380
rect 2256 4324 2312 4380
rect 2312 4324 2316 4380
rect 2252 4320 2316 4324
rect 2332 4380 2396 4384
rect 2332 4324 2336 4380
rect 2336 4324 2392 4380
rect 2392 4324 2396 4380
rect 2332 4320 2396 4324
rect 2412 4380 2476 4384
rect 2412 4324 2416 4380
rect 2416 4324 2472 4380
rect 2472 4324 2476 4380
rect 2412 4320 2476 4324
rect 2492 4380 2556 4384
rect 2492 4324 2496 4380
rect 2496 4324 2552 4380
rect 2552 4324 2556 4380
rect 2492 4320 2556 4324
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 4332 4380 4396 4384
rect 4332 4324 4336 4380
rect 4336 4324 4392 4380
rect 4392 4324 4396 4380
rect 4332 4320 4396 4324
rect 4412 4380 4476 4384
rect 4412 4324 4416 4380
rect 4416 4324 4472 4380
rect 4472 4324 4476 4380
rect 4412 4320 4476 4324
rect 4492 4380 4556 4384
rect 4492 4324 4496 4380
rect 4496 4324 4552 4380
rect 4552 4324 4556 4380
rect 4492 4320 4556 4324
rect 6252 4380 6316 4384
rect 6252 4324 6256 4380
rect 6256 4324 6312 4380
rect 6312 4324 6316 4380
rect 6252 4320 6316 4324
rect 6332 4380 6396 4384
rect 6332 4324 6336 4380
rect 6336 4324 6392 4380
rect 6392 4324 6396 4380
rect 6332 4320 6396 4324
rect 6412 4380 6476 4384
rect 6412 4324 6416 4380
rect 6416 4324 6472 4380
rect 6472 4324 6476 4380
rect 6412 4320 6476 4324
rect 6492 4380 6556 4384
rect 6492 4324 6496 4380
rect 6496 4324 6552 4380
rect 6552 4324 6556 4380
rect 6492 4320 6556 4324
rect 8252 4380 8316 4384
rect 8252 4324 8256 4380
rect 8256 4324 8312 4380
rect 8312 4324 8316 4380
rect 8252 4320 8316 4324
rect 8332 4380 8396 4384
rect 8332 4324 8336 4380
rect 8336 4324 8392 4380
rect 8392 4324 8396 4380
rect 8332 4320 8396 4324
rect 8412 4380 8476 4384
rect 8412 4324 8416 4380
rect 8416 4324 8472 4380
rect 8472 4324 8476 4380
rect 8412 4320 8476 4324
rect 8492 4380 8556 4384
rect 8492 4324 8496 4380
rect 8496 4324 8552 4380
rect 8552 4324 8556 4380
rect 8492 4320 8556 4324
rect 10252 4380 10316 4384
rect 10252 4324 10256 4380
rect 10256 4324 10312 4380
rect 10312 4324 10316 4380
rect 10252 4320 10316 4324
rect 10332 4380 10396 4384
rect 10332 4324 10336 4380
rect 10336 4324 10392 4380
rect 10392 4324 10396 4380
rect 10332 4320 10396 4324
rect 10412 4380 10476 4384
rect 10412 4324 10416 4380
rect 10416 4324 10472 4380
rect 10472 4324 10476 4380
rect 10412 4320 10476 4324
rect 10492 4380 10556 4384
rect 10492 4324 10496 4380
rect 10496 4324 10552 4380
rect 10552 4324 10556 4380
rect 10492 4320 10556 4324
rect 1552 3836 1616 3840
rect 1552 3780 1556 3836
rect 1556 3780 1612 3836
rect 1612 3780 1616 3836
rect 1552 3776 1616 3780
rect 1632 3836 1696 3840
rect 1632 3780 1636 3836
rect 1636 3780 1692 3836
rect 1692 3780 1696 3836
rect 1632 3776 1696 3780
rect 1712 3836 1776 3840
rect 1712 3780 1716 3836
rect 1716 3780 1772 3836
rect 1772 3780 1776 3836
rect 1712 3776 1776 3780
rect 1792 3836 1856 3840
rect 1792 3780 1796 3836
rect 1796 3780 1852 3836
rect 1852 3780 1856 3836
rect 1792 3776 1856 3780
rect 3552 3836 3616 3840
rect 3552 3780 3556 3836
rect 3556 3780 3612 3836
rect 3612 3780 3616 3836
rect 3552 3776 3616 3780
rect 3632 3836 3696 3840
rect 3632 3780 3636 3836
rect 3636 3780 3692 3836
rect 3692 3780 3696 3836
rect 3632 3776 3696 3780
rect 3712 3836 3776 3840
rect 3712 3780 3716 3836
rect 3716 3780 3772 3836
rect 3772 3780 3776 3836
rect 3712 3776 3776 3780
rect 3792 3836 3856 3840
rect 3792 3780 3796 3836
rect 3796 3780 3852 3836
rect 3852 3780 3856 3836
rect 3792 3776 3856 3780
rect 5552 3836 5616 3840
rect 5552 3780 5556 3836
rect 5556 3780 5612 3836
rect 5612 3780 5616 3836
rect 5552 3776 5616 3780
rect 5632 3836 5696 3840
rect 5632 3780 5636 3836
rect 5636 3780 5692 3836
rect 5692 3780 5696 3836
rect 5632 3776 5696 3780
rect 5712 3836 5776 3840
rect 5712 3780 5716 3836
rect 5716 3780 5772 3836
rect 5772 3780 5776 3836
rect 5712 3776 5776 3780
rect 5792 3836 5856 3840
rect 5792 3780 5796 3836
rect 5796 3780 5852 3836
rect 5852 3780 5856 3836
rect 5792 3776 5856 3780
rect 7552 3836 7616 3840
rect 7552 3780 7556 3836
rect 7556 3780 7612 3836
rect 7612 3780 7616 3836
rect 7552 3776 7616 3780
rect 7632 3836 7696 3840
rect 7632 3780 7636 3836
rect 7636 3780 7692 3836
rect 7692 3780 7696 3836
rect 7632 3776 7696 3780
rect 7712 3836 7776 3840
rect 7712 3780 7716 3836
rect 7716 3780 7772 3836
rect 7772 3780 7776 3836
rect 7712 3776 7776 3780
rect 7792 3836 7856 3840
rect 7792 3780 7796 3836
rect 7796 3780 7852 3836
rect 7852 3780 7856 3836
rect 7792 3776 7856 3780
rect 9552 3836 9616 3840
rect 9552 3780 9556 3836
rect 9556 3780 9612 3836
rect 9612 3780 9616 3836
rect 9552 3776 9616 3780
rect 9632 3836 9696 3840
rect 9632 3780 9636 3836
rect 9636 3780 9692 3836
rect 9692 3780 9696 3836
rect 9632 3776 9696 3780
rect 9712 3836 9776 3840
rect 9712 3780 9716 3836
rect 9716 3780 9772 3836
rect 9772 3780 9776 3836
rect 9712 3776 9776 3780
rect 9792 3836 9856 3840
rect 9792 3780 9796 3836
rect 9796 3780 9852 3836
rect 9852 3780 9856 3836
rect 9792 3776 9856 3780
rect 11552 3836 11616 3840
rect 11552 3780 11556 3836
rect 11556 3780 11612 3836
rect 11612 3780 11616 3836
rect 11552 3776 11616 3780
rect 11632 3836 11696 3840
rect 11632 3780 11636 3836
rect 11636 3780 11692 3836
rect 11692 3780 11696 3836
rect 11632 3776 11696 3780
rect 11712 3836 11776 3840
rect 11712 3780 11716 3836
rect 11716 3780 11772 3836
rect 11772 3780 11776 3836
rect 11712 3776 11776 3780
rect 11792 3836 11856 3840
rect 11792 3780 11796 3836
rect 11796 3780 11852 3836
rect 11852 3780 11856 3836
rect 11792 3776 11856 3780
rect 2252 3292 2316 3296
rect 2252 3236 2256 3292
rect 2256 3236 2312 3292
rect 2312 3236 2316 3292
rect 2252 3232 2316 3236
rect 2332 3292 2396 3296
rect 2332 3236 2336 3292
rect 2336 3236 2392 3292
rect 2392 3236 2396 3292
rect 2332 3232 2396 3236
rect 2412 3292 2476 3296
rect 2412 3236 2416 3292
rect 2416 3236 2472 3292
rect 2472 3236 2476 3292
rect 2412 3232 2476 3236
rect 2492 3292 2556 3296
rect 2492 3236 2496 3292
rect 2496 3236 2552 3292
rect 2552 3236 2556 3292
rect 2492 3232 2556 3236
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 4332 3292 4396 3296
rect 4332 3236 4336 3292
rect 4336 3236 4392 3292
rect 4392 3236 4396 3292
rect 4332 3232 4396 3236
rect 4412 3292 4476 3296
rect 4412 3236 4416 3292
rect 4416 3236 4472 3292
rect 4472 3236 4476 3292
rect 4412 3232 4476 3236
rect 4492 3292 4556 3296
rect 4492 3236 4496 3292
rect 4496 3236 4552 3292
rect 4552 3236 4556 3292
rect 4492 3232 4556 3236
rect 6252 3292 6316 3296
rect 6252 3236 6256 3292
rect 6256 3236 6312 3292
rect 6312 3236 6316 3292
rect 6252 3232 6316 3236
rect 6332 3292 6396 3296
rect 6332 3236 6336 3292
rect 6336 3236 6392 3292
rect 6392 3236 6396 3292
rect 6332 3232 6396 3236
rect 6412 3292 6476 3296
rect 6412 3236 6416 3292
rect 6416 3236 6472 3292
rect 6472 3236 6476 3292
rect 6412 3232 6476 3236
rect 6492 3292 6556 3296
rect 6492 3236 6496 3292
rect 6496 3236 6552 3292
rect 6552 3236 6556 3292
rect 6492 3232 6556 3236
rect 8252 3292 8316 3296
rect 8252 3236 8256 3292
rect 8256 3236 8312 3292
rect 8312 3236 8316 3292
rect 8252 3232 8316 3236
rect 8332 3292 8396 3296
rect 8332 3236 8336 3292
rect 8336 3236 8392 3292
rect 8392 3236 8396 3292
rect 8332 3232 8396 3236
rect 8412 3292 8476 3296
rect 8412 3236 8416 3292
rect 8416 3236 8472 3292
rect 8472 3236 8476 3292
rect 8412 3232 8476 3236
rect 8492 3292 8556 3296
rect 8492 3236 8496 3292
rect 8496 3236 8552 3292
rect 8552 3236 8556 3292
rect 8492 3232 8556 3236
rect 10252 3292 10316 3296
rect 10252 3236 10256 3292
rect 10256 3236 10312 3292
rect 10312 3236 10316 3292
rect 10252 3232 10316 3236
rect 10332 3292 10396 3296
rect 10332 3236 10336 3292
rect 10336 3236 10392 3292
rect 10392 3236 10396 3292
rect 10332 3232 10396 3236
rect 10412 3292 10476 3296
rect 10412 3236 10416 3292
rect 10416 3236 10472 3292
rect 10472 3236 10476 3292
rect 10412 3232 10476 3236
rect 10492 3292 10556 3296
rect 10492 3236 10496 3292
rect 10496 3236 10552 3292
rect 10552 3236 10556 3292
rect 10492 3232 10556 3236
rect 1552 2748 1616 2752
rect 1552 2692 1556 2748
rect 1556 2692 1612 2748
rect 1612 2692 1616 2748
rect 1552 2688 1616 2692
rect 1632 2748 1696 2752
rect 1632 2692 1636 2748
rect 1636 2692 1692 2748
rect 1692 2692 1696 2748
rect 1632 2688 1696 2692
rect 1712 2748 1776 2752
rect 1712 2692 1716 2748
rect 1716 2692 1772 2748
rect 1772 2692 1776 2748
rect 1712 2688 1776 2692
rect 1792 2748 1856 2752
rect 1792 2692 1796 2748
rect 1796 2692 1852 2748
rect 1852 2692 1856 2748
rect 1792 2688 1856 2692
rect 3552 2748 3616 2752
rect 3552 2692 3556 2748
rect 3556 2692 3612 2748
rect 3612 2692 3616 2748
rect 3552 2688 3616 2692
rect 3632 2748 3696 2752
rect 3632 2692 3636 2748
rect 3636 2692 3692 2748
rect 3692 2692 3696 2748
rect 3632 2688 3696 2692
rect 3712 2748 3776 2752
rect 3712 2692 3716 2748
rect 3716 2692 3772 2748
rect 3772 2692 3776 2748
rect 3712 2688 3776 2692
rect 3792 2748 3856 2752
rect 3792 2692 3796 2748
rect 3796 2692 3852 2748
rect 3852 2692 3856 2748
rect 3792 2688 3856 2692
rect 5552 2748 5616 2752
rect 5552 2692 5556 2748
rect 5556 2692 5612 2748
rect 5612 2692 5616 2748
rect 5552 2688 5616 2692
rect 5632 2748 5696 2752
rect 5632 2692 5636 2748
rect 5636 2692 5692 2748
rect 5692 2692 5696 2748
rect 5632 2688 5696 2692
rect 5712 2748 5776 2752
rect 5712 2692 5716 2748
rect 5716 2692 5772 2748
rect 5772 2692 5776 2748
rect 5712 2688 5776 2692
rect 5792 2748 5856 2752
rect 5792 2692 5796 2748
rect 5796 2692 5852 2748
rect 5852 2692 5856 2748
rect 5792 2688 5856 2692
rect 7552 2748 7616 2752
rect 7552 2692 7556 2748
rect 7556 2692 7612 2748
rect 7612 2692 7616 2748
rect 7552 2688 7616 2692
rect 7632 2748 7696 2752
rect 7632 2692 7636 2748
rect 7636 2692 7692 2748
rect 7692 2692 7696 2748
rect 7632 2688 7696 2692
rect 7712 2748 7776 2752
rect 7712 2692 7716 2748
rect 7716 2692 7772 2748
rect 7772 2692 7776 2748
rect 7712 2688 7776 2692
rect 7792 2748 7856 2752
rect 7792 2692 7796 2748
rect 7796 2692 7852 2748
rect 7852 2692 7856 2748
rect 7792 2688 7856 2692
rect 9552 2748 9616 2752
rect 9552 2692 9556 2748
rect 9556 2692 9612 2748
rect 9612 2692 9616 2748
rect 9552 2688 9616 2692
rect 9632 2748 9696 2752
rect 9632 2692 9636 2748
rect 9636 2692 9692 2748
rect 9692 2692 9696 2748
rect 9632 2688 9696 2692
rect 9712 2748 9776 2752
rect 9712 2692 9716 2748
rect 9716 2692 9772 2748
rect 9772 2692 9776 2748
rect 9712 2688 9776 2692
rect 9792 2748 9856 2752
rect 9792 2692 9796 2748
rect 9796 2692 9852 2748
rect 9852 2692 9856 2748
rect 9792 2688 9856 2692
rect 11552 2748 11616 2752
rect 11552 2692 11556 2748
rect 11556 2692 11612 2748
rect 11612 2692 11616 2748
rect 11552 2688 11616 2692
rect 11632 2748 11696 2752
rect 11632 2692 11636 2748
rect 11636 2692 11692 2748
rect 11692 2692 11696 2748
rect 11632 2688 11696 2692
rect 11712 2748 11776 2752
rect 11712 2692 11716 2748
rect 11716 2692 11772 2748
rect 11772 2692 11776 2748
rect 11712 2688 11776 2692
rect 11792 2748 11856 2752
rect 11792 2692 11796 2748
rect 11796 2692 11852 2748
rect 11852 2692 11856 2748
rect 11792 2688 11856 2692
rect 2252 2204 2316 2208
rect 2252 2148 2256 2204
rect 2256 2148 2312 2204
rect 2312 2148 2316 2204
rect 2252 2144 2316 2148
rect 2332 2204 2396 2208
rect 2332 2148 2336 2204
rect 2336 2148 2392 2204
rect 2392 2148 2396 2204
rect 2332 2144 2396 2148
rect 2412 2204 2476 2208
rect 2412 2148 2416 2204
rect 2416 2148 2472 2204
rect 2472 2148 2476 2204
rect 2412 2144 2476 2148
rect 2492 2204 2556 2208
rect 2492 2148 2496 2204
rect 2496 2148 2552 2204
rect 2552 2148 2556 2204
rect 2492 2144 2556 2148
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 4332 2204 4396 2208
rect 4332 2148 4336 2204
rect 4336 2148 4392 2204
rect 4392 2148 4396 2204
rect 4332 2144 4396 2148
rect 4412 2204 4476 2208
rect 4412 2148 4416 2204
rect 4416 2148 4472 2204
rect 4472 2148 4476 2204
rect 4412 2144 4476 2148
rect 4492 2204 4556 2208
rect 4492 2148 4496 2204
rect 4496 2148 4552 2204
rect 4552 2148 4556 2204
rect 4492 2144 4556 2148
rect 6252 2204 6316 2208
rect 6252 2148 6256 2204
rect 6256 2148 6312 2204
rect 6312 2148 6316 2204
rect 6252 2144 6316 2148
rect 6332 2204 6396 2208
rect 6332 2148 6336 2204
rect 6336 2148 6392 2204
rect 6392 2148 6396 2204
rect 6332 2144 6396 2148
rect 6412 2204 6476 2208
rect 6412 2148 6416 2204
rect 6416 2148 6472 2204
rect 6472 2148 6476 2204
rect 6412 2144 6476 2148
rect 6492 2204 6556 2208
rect 6492 2148 6496 2204
rect 6496 2148 6552 2204
rect 6552 2148 6556 2204
rect 6492 2144 6556 2148
rect 8252 2204 8316 2208
rect 8252 2148 8256 2204
rect 8256 2148 8312 2204
rect 8312 2148 8316 2204
rect 8252 2144 8316 2148
rect 8332 2204 8396 2208
rect 8332 2148 8336 2204
rect 8336 2148 8392 2204
rect 8392 2148 8396 2204
rect 8332 2144 8396 2148
rect 8412 2204 8476 2208
rect 8412 2148 8416 2204
rect 8416 2148 8472 2204
rect 8472 2148 8476 2204
rect 8412 2144 8476 2148
rect 8492 2204 8556 2208
rect 8492 2148 8496 2204
rect 8496 2148 8552 2204
rect 8552 2148 8556 2204
rect 8492 2144 8556 2148
rect 10252 2204 10316 2208
rect 10252 2148 10256 2204
rect 10256 2148 10312 2204
rect 10312 2148 10316 2204
rect 10252 2144 10316 2148
rect 10332 2204 10396 2208
rect 10332 2148 10336 2204
rect 10336 2148 10392 2204
rect 10392 2148 10396 2204
rect 10332 2144 10396 2148
rect 10412 2204 10476 2208
rect 10412 2148 10416 2204
rect 10416 2148 10472 2204
rect 10472 2148 10476 2204
rect 10412 2144 10476 2148
rect 10492 2204 10556 2208
rect 10492 2148 10496 2204
rect 10496 2148 10552 2204
rect 10552 2148 10556 2204
rect 10492 2144 10556 2148
<< metal4 >>
rect -1076 15194 -756 15236
rect -1076 14958 -1034 15194
rect -798 14958 -756 15194
rect -1076 11594 -756 14958
rect -1076 11358 -1034 11594
rect -798 11358 -756 11594
rect -1076 9594 -756 11358
rect -1076 9358 -1034 9594
rect -798 9358 -756 9594
rect -1076 7594 -756 9358
rect -1076 7358 -1034 7594
rect -798 7358 -756 7594
rect -1076 5594 -756 7358
rect -1076 5358 -1034 5594
rect -798 5358 -756 5594
rect -1076 3594 -756 5358
rect -1076 3358 -1034 3594
rect -798 3358 -756 3594
rect -1076 274 -756 3358
rect -416 14534 -96 14576
rect -416 14298 -374 14534
rect -138 14298 -96 14534
rect -416 12894 -96 14298
rect -416 12658 -374 12894
rect -138 12658 -96 12894
rect -416 10894 -96 12658
rect -416 10658 -374 10894
rect -138 10658 -96 10894
rect -416 8894 -96 10658
rect -416 8658 -374 8894
rect -138 8658 -96 8894
rect -416 6894 -96 8658
rect -416 6658 -374 6894
rect -138 6658 -96 6894
rect -416 4894 -96 6658
rect -416 4658 -374 4894
rect -138 4658 -96 4894
rect -416 2894 -96 4658
rect -416 2658 -374 2894
rect -138 2658 -96 2894
rect -416 934 -96 2658
rect -416 698 -374 934
rect -138 698 -96 934
rect -416 656 -96 698
rect 1524 14534 1884 15236
rect 1524 14298 1586 14534
rect 1822 14298 1884 14534
rect 1524 12894 1884 14298
rect 1524 12658 1586 12894
rect 1822 12658 1884 12894
rect 1524 12544 1884 12658
rect 1524 12480 1552 12544
rect 1616 12480 1632 12544
rect 1696 12480 1712 12544
rect 1776 12480 1792 12544
rect 1856 12480 1884 12544
rect 1524 11456 1884 12480
rect 1524 11392 1552 11456
rect 1616 11392 1632 11456
rect 1696 11392 1712 11456
rect 1776 11392 1792 11456
rect 1856 11392 1884 11456
rect 1524 10894 1884 11392
rect 1524 10658 1586 10894
rect 1822 10658 1884 10894
rect 1524 10368 1884 10658
rect 1524 10304 1552 10368
rect 1616 10304 1632 10368
rect 1696 10304 1712 10368
rect 1776 10304 1792 10368
rect 1856 10304 1884 10368
rect 1524 9280 1884 10304
rect 1524 9216 1552 9280
rect 1616 9216 1632 9280
rect 1696 9216 1712 9280
rect 1776 9216 1792 9280
rect 1856 9216 1884 9280
rect 1524 8894 1884 9216
rect 1524 8658 1586 8894
rect 1822 8658 1884 8894
rect 1524 8192 1884 8658
rect 1524 8128 1552 8192
rect 1616 8128 1632 8192
rect 1696 8128 1712 8192
rect 1776 8128 1792 8192
rect 1856 8128 1884 8192
rect 1524 7104 1884 8128
rect 1524 7040 1552 7104
rect 1616 7040 1632 7104
rect 1696 7040 1712 7104
rect 1776 7040 1792 7104
rect 1856 7040 1884 7104
rect 1524 6894 1884 7040
rect 1524 6658 1586 6894
rect 1822 6658 1884 6894
rect 1524 6016 1884 6658
rect 1524 5952 1552 6016
rect 1616 5952 1632 6016
rect 1696 5952 1712 6016
rect 1776 5952 1792 6016
rect 1856 5952 1884 6016
rect 1524 4928 1884 5952
rect 1524 4864 1552 4928
rect 1616 4894 1632 4928
rect 1696 4894 1712 4928
rect 1776 4894 1792 4928
rect 1856 4864 1884 4928
rect 1524 4658 1586 4864
rect 1822 4658 1884 4864
rect 1524 3840 1884 4658
rect 1524 3776 1552 3840
rect 1616 3776 1632 3840
rect 1696 3776 1712 3840
rect 1776 3776 1792 3840
rect 1856 3776 1884 3840
rect 1524 2894 1884 3776
rect 1524 2752 1586 2894
rect 1822 2752 1884 2894
rect 1524 2688 1552 2752
rect 1856 2688 1884 2752
rect 1524 2658 1586 2688
rect 1822 2658 1884 2688
rect 1524 934 1884 2658
rect 1524 698 1586 934
rect 1822 698 1884 934
rect -1076 38 -1034 274
rect -798 38 -756 274
rect -1076 -4 -756 38
rect 1524 -4 1884 698
rect 2224 15194 2584 15236
rect 2224 14958 2286 15194
rect 2522 14958 2584 15194
rect 2224 13088 2584 14958
rect 2224 13024 2252 13088
rect 2316 13024 2332 13088
rect 2396 13024 2412 13088
rect 2476 13024 2492 13088
rect 2556 13024 2584 13088
rect 2224 12000 2584 13024
rect 2224 11936 2252 12000
rect 2316 11936 2332 12000
rect 2396 11936 2412 12000
rect 2476 11936 2492 12000
rect 2556 11936 2584 12000
rect 2224 11594 2584 11936
rect 2224 11358 2286 11594
rect 2522 11358 2584 11594
rect 2224 10912 2584 11358
rect 2224 10848 2252 10912
rect 2316 10848 2332 10912
rect 2396 10848 2412 10912
rect 2476 10848 2492 10912
rect 2556 10848 2584 10912
rect 2224 9824 2584 10848
rect 2224 9760 2252 9824
rect 2316 9760 2332 9824
rect 2396 9760 2412 9824
rect 2476 9760 2492 9824
rect 2556 9760 2584 9824
rect 2224 9594 2584 9760
rect 2224 9358 2286 9594
rect 2522 9358 2584 9594
rect 2224 8736 2584 9358
rect 2224 8672 2252 8736
rect 2316 8672 2332 8736
rect 2396 8672 2412 8736
rect 2476 8672 2492 8736
rect 2556 8672 2584 8736
rect 2224 7648 2584 8672
rect 2224 7584 2252 7648
rect 2316 7594 2332 7648
rect 2396 7594 2412 7648
rect 2476 7594 2492 7648
rect 2556 7584 2584 7648
rect 2224 7358 2286 7584
rect 2522 7358 2584 7584
rect 2224 6560 2584 7358
rect 2224 6496 2252 6560
rect 2316 6496 2332 6560
rect 2396 6496 2412 6560
rect 2476 6496 2492 6560
rect 2556 6496 2584 6560
rect 2224 5594 2584 6496
rect 2224 5472 2286 5594
rect 2522 5472 2584 5594
rect 2224 5408 2252 5472
rect 2556 5408 2584 5472
rect 2224 5358 2286 5408
rect 2522 5358 2584 5408
rect 2224 4384 2584 5358
rect 2224 4320 2252 4384
rect 2316 4320 2332 4384
rect 2396 4320 2412 4384
rect 2476 4320 2492 4384
rect 2556 4320 2584 4384
rect 2224 3594 2584 4320
rect 2224 3358 2286 3594
rect 2522 3358 2584 3594
rect 2224 3296 2584 3358
rect 2224 3232 2252 3296
rect 2316 3232 2332 3296
rect 2396 3232 2412 3296
rect 2476 3232 2492 3296
rect 2556 3232 2584 3296
rect 2224 2208 2584 3232
rect 2224 2144 2252 2208
rect 2316 2144 2332 2208
rect 2396 2144 2412 2208
rect 2476 2144 2492 2208
rect 2556 2144 2584 2208
rect 2224 274 2584 2144
rect 2224 38 2286 274
rect 2522 38 2584 274
rect 2224 -4 2584 38
rect 3524 14534 3884 15236
rect 3524 14298 3586 14534
rect 3822 14298 3884 14534
rect 3524 12894 3884 14298
rect 3524 12658 3586 12894
rect 3822 12658 3884 12894
rect 3524 12544 3884 12658
rect 3524 12480 3552 12544
rect 3616 12480 3632 12544
rect 3696 12480 3712 12544
rect 3776 12480 3792 12544
rect 3856 12480 3884 12544
rect 3524 11456 3884 12480
rect 3524 11392 3552 11456
rect 3616 11392 3632 11456
rect 3696 11392 3712 11456
rect 3776 11392 3792 11456
rect 3856 11392 3884 11456
rect 3524 10894 3884 11392
rect 3524 10658 3586 10894
rect 3822 10658 3884 10894
rect 3524 10368 3884 10658
rect 3524 10304 3552 10368
rect 3616 10304 3632 10368
rect 3696 10304 3712 10368
rect 3776 10304 3792 10368
rect 3856 10304 3884 10368
rect 3524 9280 3884 10304
rect 3524 9216 3552 9280
rect 3616 9216 3632 9280
rect 3696 9216 3712 9280
rect 3776 9216 3792 9280
rect 3856 9216 3884 9280
rect 3524 8894 3884 9216
rect 3524 8658 3586 8894
rect 3822 8658 3884 8894
rect 3524 8192 3884 8658
rect 3524 8128 3552 8192
rect 3616 8128 3632 8192
rect 3696 8128 3712 8192
rect 3776 8128 3792 8192
rect 3856 8128 3884 8192
rect 3524 7104 3884 8128
rect 3524 7040 3552 7104
rect 3616 7040 3632 7104
rect 3696 7040 3712 7104
rect 3776 7040 3792 7104
rect 3856 7040 3884 7104
rect 3524 6894 3884 7040
rect 3524 6658 3586 6894
rect 3822 6658 3884 6894
rect 3524 6016 3884 6658
rect 3524 5952 3552 6016
rect 3616 5952 3632 6016
rect 3696 5952 3712 6016
rect 3776 5952 3792 6016
rect 3856 5952 3884 6016
rect 3524 4928 3884 5952
rect 3524 4864 3552 4928
rect 3616 4894 3632 4928
rect 3696 4894 3712 4928
rect 3776 4894 3792 4928
rect 3856 4864 3884 4928
rect 3524 4658 3586 4864
rect 3822 4658 3884 4864
rect 3524 3840 3884 4658
rect 3524 3776 3552 3840
rect 3616 3776 3632 3840
rect 3696 3776 3712 3840
rect 3776 3776 3792 3840
rect 3856 3776 3884 3840
rect 3524 2894 3884 3776
rect 3524 2752 3586 2894
rect 3822 2752 3884 2894
rect 3524 2688 3552 2752
rect 3856 2688 3884 2752
rect 3524 2658 3586 2688
rect 3822 2658 3884 2688
rect 3524 934 3884 2658
rect 3524 698 3586 934
rect 3822 698 3884 934
rect 3524 -4 3884 698
rect 4224 15194 4584 15236
rect 4224 14958 4286 15194
rect 4522 14958 4584 15194
rect 4224 13088 4584 14958
rect 4224 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4584 13088
rect 4224 12000 4584 13024
rect 4224 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4584 12000
rect 4224 11594 4584 11936
rect 4224 11358 4286 11594
rect 4522 11358 4584 11594
rect 4224 10912 4584 11358
rect 4224 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4584 10912
rect 4224 9824 4584 10848
rect 4224 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4584 9824
rect 4224 9594 4584 9760
rect 4224 9358 4286 9594
rect 4522 9358 4584 9594
rect 4224 8736 4584 9358
rect 4224 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4584 8736
rect 4224 7648 4584 8672
rect 4224 7584 4252 7648
rect 4316 7594 4332 7648
rect 4396 7594 4412 7648
rect 4476 7594 4492 7648
rect 4556 7584 4584 7648
rect 4224 7358 4286 7584
rect 4522 7358 4584 7584
rect 4224 6560 4584 7358
rect 4224 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4584 6560
rect 4224 5594 4584 6496
rect 4224 5472 4286 5594
rect 4522 5472 4584 5594
rect 4224 5408 4252 5472
rect 4556 5408 4584 5472
rect 4224 5358 4286 5408
rect 4522 5358 4584 5408
rect 4224 4384 4584 5358
rect 4224 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4584 4384
rect 4224 3594 4584 4320
rect 4224 3358 4286 3594
rect 4522 3358 4584 3594
rect 4224 3296 4584 3358
rect 4224 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4584 3296
rect 4224 2208 4584 3232
rect 4224 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4584 2208
rect 4224 274 4584 2144
rect 4224 38 4286 274
rect 4522 38 4584 274
rect 4224 -4 4584 38
rect 5524 14534 5884 15236
rect 5524 14298 5586 14534
rect 5822 14298 5884 14534
rect 5524 12894 5884 14298
rect 5524 12658 5586 12894
rect 5822 12658 5884 12894
rect 5524 12544 5884 12658
rect 5524 12480 5552 12544
rect 5616 12480 5632 12544
rect 5696 12480 5712 12544
rect 5776 12480 5792 12544
rect 5856 12480 5884 12544
rect 5524 11456 5884 12480
rect 5524 11392 5552 11456
rect 5616 11392 5632 11456
rect 5696 11392 5712 11456
rect 5776 11392 5792 11456
rect 5856 11392 5884 11456
rect 5524 10894 5884 11392
rect 5524 10658 5586 10894
rect 5822 10658 5884 10894
rect 5524 10368 5884 10658
rect 5524 10304 5552 10368
rect 5616 10304 5632 10368
rect 5696 10304 5712 10368
rect 5776 10304 5792 10368
rect 5856 10304 5884 10368
rect 5524 9280 5884 10304
rect 5524 9216 5552 9280
rect 5616 9216 5632 9280
rect 5696 9216 5712 9280
rect 5776 9216 5792 9280
rect 5856 9216 5884 9280
rect 5524 8894 5884 9216
rect 5524 8658 5586 8894
rect 5822 8658 5884 8894
rect 5524 8192 5884 8658
rect 5524 8128 5552 8192
rect 5616 8128 5632 8192
rect 5696 8128 5712 8192
rect 5776 8128 5792 8192
rect 5856 8128 5884 8192
rect 5524 7104 5884 8128
rect 5524 7040 5552 7104
rect 5616 7040 5632 7104
rect 5696 7040 5712 7104
rect 5776 7040 5792 7104
rect 5856 7040 5884 7104
rect 5524 6894 5884 7040
rect 5524 6658 5586 6894
rect 5822 6658 5884 6894
rect 5524 6016 5884 6658
rect 5524 5952 5552 6016
rect 5616 5952 5632 6016
rect 5696 5952 5712 6016
rect 5776 5952 5792 6016
rect 5856 5952 5884 6016
rect 5524 4928 5884 5952
rect 5524 4864 5552 4928
rect 5616 4894 5632 4928
rect 5696 4894 5712 4928
rect 5776 4894 5792 4928
rect 5856 4864 5884 4928
rect 5524 4658 5586 4864
rect 5822 4658 5884 4864
rect 5524 3840 5884 4658
rect 5524 3776 5552 3840
rect 5616 3776 5632 3840
rect 5696 3776 5712 3840
rect 5776 3776 5792 3840
rect 5856 3776 5884 3840
rect 5524 2894 5884 3776
rect 5524 2752 5586 2894
rect 5822 2752 5884 2894
rect 5524 2688 5552 2752
rect 5856 2688 5884 2752
rect 5524 2658 5586 2688
rect 5822 2658 5884 2688
rect 5524 934 5884 2658
rect 5524 698 5586 934
rect 5822 698 5884 934
rect 5524 -4 5884 698
rect 6224 15194 6584 15236
rect 6224 14958 6286 15194
rect 6522 14958 6584 15194
rect 6224 13088 6584 14958
rect 6224 13024 6252 13088
rect 6316 13024 6332 13088
rect 6396 13024 6412 13088
rect 6476 13024 6492 13088
rect 6556 13024 6584 13088
rect 6224 12000 6584 13024
rect 6224 11936 6252 12000
rect 6316 11936 6332 12000
rect 6396 11936 6412 12000
rect 6476 11936 6492 12000
rect 6556 11936 6584 12000
rect 6224 11594 6584 11936
rect 6224 11358 6286 11594
rect 6522 11358 6584 11594
rect 6224 10912 6584 11358
rect 6224 10848 6252 10912
rect 6316 10848 6332 10912
rect 6396 10848 6412 10912
rect 6476 10848 6492 10912
rect 6556 10848 6584 10912
rect 6224 9824 6584 10848
rect 6224 9760 6252 9824
rect 6316 9760 6332 9824
rect 6396 9760 6412 9824
rect 6476 9760 6492 9824
rect 6556 9760 6584 9824
rect 6224 9594 6584 9760
rect 6224 9358 6286 9594
rect 6522 9358 6584 9594
rect 6224 8736 6584 9358
rect 6224 8672 6252 8736
rect 6316 8672 6332 8736
rect 6396 8672 6412 8736
rect 6476 8672 6492 8736
rect 6556 8672 6584 8736
rect 6224 7648 6584 8672
rect 6224 7584 6252 7648
rect 6316 7594 6332 7648
rect 6396 7594 6412 7648
rect 6476 7594 6492 7648
rect 6556 7584 6584 7648
rect 6224 7358 6286 7584
rect 6522 7358 6584 7584
rect 6224 6560 6584 7358
rect 6224 6496 6252 6560
rect 6316 6496 6332 6560
rect 6396 6496 6412 6560
rect 6476 6496 6492 6560
rect 6556 6496 6584 6560
rect 6224 5594 6584 6496
rect 6224 5472 6286 5594
rect 6522 5472 6584 5594
rect 6224 5408 6252 5472
rect 6556 5408 6584 5472
rect 6224 5358 6286 5408
rect 6522 5358 6584 5408
rect 6224 4384 6584 5358
rect 6224 4320 6252 4384
rect 6316 4320 6332 4384
rect 6396 4320 6412 4384
rect 6476 4320 6492 4384
rect 6556 4320 6584 4384
rect 6224 3594 6584 4320
rect 6224 3358 6286 3594
rect 6522 3358 6584 3594
rect 6224 3296 6584 3358
rect 6224 3232 6252 3296
rect 6316 3232 6332 3296
rect 6396 3232 6412 3296
rect 6476 3232 6492 3296
rect 6556 3232 6584 3296
rect 6224 2208 6584 3232
rect 6224 2144 6252 2208
rect 6316 2144 6332 2208
rect 6396 2144 6412 2208
rect 6476 2144 6492 2208
rect 6556 2144 6584 2208
rect 6224 274 6584 2144
rect 6224 38 6286 274
rect 6522 38 6584 274
rect 6224 -4 6584 38
rect 7524 14534 7884 15236
rect 7524 14298 7586 14534
rect 7822 14298 7884 14534
rect 7524 12894 7884 14298
rect 7524 12658 7586 12894
rect 7822 12658 7884 12894
rect 7524 12544 7884 12658
rect 7524 12480 7552 12544
rect 7616 12480 7632 12544
rect 7696 12480 7712 12544
rect 7776 12480 7792 12544
rect 7856 12480 7884 12544
rect 7524 11456 7884 12480
rect 7524 11392 7552 11456
rect 7616 11392 7632 11456
rect 7696 11392 7712 11456
rect 7776 11392 7792 11456
rect 7856 11392 7884 11456
rect 7524 10894 7884 11392
rect 7524 10658 7586 10894
rect 7822 10658 7884 10894
rect 7524 10368 7884 10658
rect 7524 10304 7552 10368
rect 7616 10304 7632 10368
rect 7696 10304 7712 10368
rect 7776 10304 7792 10368
rect 7856 10304 7884 10368
rect 7524 9280 7884 10304
rect 7524 9216 7552 9280
rect 7616 9216 7632 9280
rect 7696 9216 7712 9280
rect 7776 9216 7792 9280
rect 7856 9216 7884 9280
rect 7524 8894 7884 9216
rect 7524 8658 7586 8894
rect 7822 8658 7884 8894
rect 7524 8192 7884 8658
rect 7524 8128 7552 8192
rect 7616 8128 7632 8192
rect 7696 8128 7712 8192
rect 7776 8128 7792 8192
rect 7856 8128 7884 8192
rect 7524 7104 7884 8128
rect 7524 7040 7552 7104
rect 7616 7040 7632 7104
rect 7696 7040 7712 7104
rect 7776 7040 7792 7104
rect 7856 7040 7884 7104
rect 7524 6894 7884 7040
rect 7524 6658 7586 6894
rect 7822 6658 7884 6894
rect 7524 6016 7884 6658
rect 7524 5952 7552 6016
rect 7616 5952 7632 6016
rect 7696 5952 7712 6016
rect 7776 5952 7792 6016
rect 7856 5952 7884 6016
rect 7524 4928 7884 5952
rect 7524 4864 7552 4928
rect 7616 4894 7632 4928
rect 7696 4894 7712 4928
rect 7776 4894 7792 4928
rect 7856 4864 7884 4928
rect 7524 4658 7586 4864
rect 7822 4658 7884 4864
rect 7524 3840 7884 4658
rect 7524 3776 7552 3840
rect 7616 3776 7632 3840
rect 7696 3776 7712 3840
rect 7776 3776 7792 3840
rect 7856 3776 7884 3840
rect 7524 2894 7884 3776
rect 7524 2752 7586 2894
rect 7822 2752 7884 2894
rect 7524 2688 7552 2752
rect 7856 2688 7884 2752
rect 7524 2658 7586 2688
rect 7822 2658 7884 2688
rect 7524 934 7884 2658
rect 7524 698 7586 934
rect 7822 698 7884 934
rect 7524 -4 7884 698
rect 8224 15194 8584 15236
rect 8224 14958 8286 15194
rect 8522 14958 8584 15194
rect 8224 13088 8584 14958
rect 8224 13024 8252 13088
rect 8316 13024 8332 13088
rect 8396 13024 8412 13088
rect 8476 13024 8492 13088
rect 8556 13024 8584 13088
rect 8224 12000 8584 13024
rect 8224 11936 8252 12000
rect 8316 11936 8332 12000
rect 8396 11936 8412 12000
rect 8476 11936 8492 12000
rect 8556 11936 8584 12000
rect 8224 11594 8584 11936
rect 8224 11358 8286 11594
rect 8522 11358 8584 11594
rect 8224 10912 8584 11358
rect 8224 10848 8252 10912
rect 8316 10848 8332 10912
rect 8396 10848 8412 10912
rect 8476 10848 8492 10912
rect 8556 10848 8584 10912
rect 8224 9824 8584 10848
rect 8224 9760 8252 9824
rect 8316 9760 8332 9824
rect 8396 9760 8412 9824
rect 8476 9760 8492 9824
rect 8556 9760 8584 9824
rect 8224 9594 8584 9760
rect 8224 9358 8286 9594
rect 8522 9358 8584 9594
rect 8224 8736 8584 9358
rect 8224 8672 8252 8736
rect 8316 8672 8332 8736
rect 8396 8672 8412 8736
rect 8476 8672 8492 8736
rect 8556 8672 8584 8736
rect 8224 7648 8584 8672
rect 8224 7584 8252 7648
rect 8316 7594 8332 7648
rect 8396 7594 8412 7648
rect 8476 7594 8492 7648
rect 8556 7584 8584 7648
rect 8224 7358 8286 7584
rect 8522 7358 8584 7584
rect 8224 6560 8584 7358
rect 8224 6496 8252 6560
rect 8316 6496 8332 6560
rect 8396 6496 8412 6560
rect 8476 6496 8492 6560
rect 8556 6496 8584 6560
rect 8224 5594 8584 6496
rect 8224 5472 8286 5594
rect 8522 5472 8584 5594
rect 8224 5408 8252 5472
rect 8556 5408 8584 5472
rect 8224 5358 8286 5408
rect 8522 5358 8584 5408
rect 8224 4384 8584 5358
rect 8224 4320 8252 4384
rect 8316 4320 8332 4384
rect 8396 4320 8412 4384
rect 8476 4320 8492 4384
rect 8556 4320 8584 4384
rect 8224 3594 8584 4320
rect 8224 3358 8286 3594
rect 8522 3358 8584 3594
rect 8224 3296 8584 3358
rect 8224 3232 8252 3296
rect 8316 3232 8332 3296
rect 8396 3232 8412 3296
rect 8476 3232 8492 3296
rect 8556 3232 8584 3296
rect 8224 2208 8584 3232
rect 8224 2144 8252 2208
rect 8316 2144 8332 2208
rect 8396 2144 8412 2208
rect 8476 2144 8492 2208
rect 8556 2144 8584 2208
rect 8224 274 8584 2144
rect 8224 38 8286 274
rect 8522 38 8584 274
rect 8224 -4 8584 38
rect 9524 14534 9884 15236
rect 9524 14298 9586 14534
rect 9822 14298 9884 14534
rect 9524 12894 9884 14298
rect 9524 12658 9586 12894
rect 9822 12658 9884 12894
rect 9524 12544 9884 12658
rect 9524 12480 9552 12544
rect 9616 12480 9632 12544
rect 9696 12480 9712 12544
rect 9776 12480 9792 12544
rect 9856 12480 9884 12544
rect 9524 11456 9884 12480
rect 9524 11392 9552 11456
rect 9616 11392 9632 11456
rect 9696 11392 9712 11456
rect 9776 11392 9792 11456
rect 9856 11392 9884 11456
rect 9524 10894 9884 11392
rect 9524 10658 9586 10894
rect 9822 10658 9884 10894
rect 9524 10368 9884 10658
rect 9524 10304 9552 10368
rect 9616 10304 9632 10368
rect 9696 10304 9712 10368
rect 9776 10304 9792 10368
rect 9856 10304 9884 10368
rect 9524 9280 9884 10304
rect 9524 9216 9552 9280
rect 9616 9216 9632 9280
rect 9696 9216 9712 9280
rect 9776 9216 9792 9280
rect 9856 9216 9884 9280
rect 9524 8894 9884 9216
rect 9524 8658 9586 8894
rect 9822 8658 9884 8894
rect 9524 8192 9884 8658
rect 9524 8128 9552 8192
rect 9616 8128 9632 8192
rect 9696 8128 9712 8192
rect 9776 8128 9792 8192
rect 9856 8128 9884 8192
rect 9524 7104 9884 8128
rect 9524 7040 9552 7104
rect 9616 7040 9632 7104
rect 9696 7040 9712 7104
rect 9776 7040 9792 7104
rect 9856 7040 9884 7104
rect 9524 6894 9884 7040
rect 9524 6658 9586 6894
rect 9822 6658 9884 6894
rect 9524 6016 9884 6658
rect 9524 5952 9552 6016
rect 9616 5952 9632 6016
rect 9696 5952 9712 6016
rect 9776 5952 9792 6016
rect 9856 5952 9884 6016
rect 9524 4928 9884 5952
rect 9524 4864 9552 4928
rect 9616 4894 9632 4928
rect 9696 4894 9712 4928
rect 9776 4894 9792 4928
rect 9856 4864 9884 4928
rect 9524 4658 9586 4864
rect 9822 4658 9884 4864
rect 9524 3840 9884 4658
rect 9524 3776 9552 3840
rect 9616 3776 9632 3840
rect 9696 3776 9712 3840
rect 9776 3776 9792 3840
rect 9856 3776 9884 3840
rect 9524 2894 9884 3776
rect 9524 2752 9586 2894
rect 9822 2752 9884 2894
rect 9524 2688 9552 2752
rect 9856 2688 9884 2752
rect 9524 2658 9586 2688
rect 9822 2658 9884 2688
rect 9524 934 9884 2658
rect 9524 698 9586 934
rect 9822 698 9884 934
rect 9524 -4 9884 698
rect 10224 15194 10584 15236
rect 10224 14958 10286 15194
rect 10522 14958 10584 15194
rect 10224 13088 10584 14958
rect 10224 13024 10252 13088
rect 10316 13024 10332 13088
rect 10396 13024 10412 13088
rect 10476 13024 10492 13088
rect 10556 13024 10584 13088
rect 10224 12000 10584 13024
rect 10224 11936 10252 12000
rect 10316 11936 10332 12000
rect 10396 11936 10412 12000
rect 10476 11936 10492 12000
rect 10556 11936 10584 12000
rect 10224 11594 10584 11936
rect 10224 11358 10286 11594
rect 10522 11358 10584 11594
rect 10224 10912 10584 11358
rect 10224 10848 10252 10912
rect 10316 10848 10332 10912
rect 10396 10848 10412 10912
rect 10476 10848 10492 10912
rect 10556 10848 10584 10912
rect 10224 9824 10584 10848
rect 10224 9760 10252 9824
rect 10316 9760 10332 9824
rect 10396 9760 10412 9824
rect 10476 9760 10492 9824
rect 10556 9760 10584 9824
rect 10224 9594 10584 9760
rect 10224 9358 10286 9594
rect 10522 9358 10584 9594
rect 10224 8736 10584 9358
rect 10224 8672 10252 8736
rect 10316 8672 10332 8736
rect 10396 8672 10412 8736
rect 10476 8672 10492 8736
rect 10556 8672 10584 8736
rect 10224 7648 10584 8672
rect 10224 7584 10252 7648
rect 10316 7594 10332 7648
rect 10396 7594 10412 7648
rect 10476 7594 10492 7648
rect 10556 7584 10584 7648
rect 10224 7358 10286 7584
rect 10522 7358 10584 7584
rect 10224 6560 10584 7358
rect 10224 6496 10252 6560
rect 10316 6496 10332 6560
rect 10396 6496 10412 6560
rect 10476 6496 10492 6560
rect 10556 6496 10584 6560
rect 10224 5594 10584 6496
rect 10224 5472 10286 5594
rect 10522 5472 10584 5594
rect 10224 5408 10252 5472
rect 10556 5408 10584 5472
rect 10224 5358 10286 5408
rect 10522 5358 10584 5408
rect 10224 4384 10584 5358
rect 10224 4320 10252 4384
rect 10316 4320 10332 4384
rect 10396 4320 10412 4384
rect 10476 4320 10492 4384
rect 10556 4320 10584 4384
rect 10224 3594 10584 4320
rect 10224 3358 10286 3594
rect 10522 3358 10584 3594
rect 10224 3296 10584 3358
rect 10224 3232 10252 3296
rect 10316 3232 10332 3296
rect 10396 3232 10412 3296
rect 10476 3232 10492 3296
rect 10556 3232 10584 3296
rect 10224 2208 10584 3232
rect 10224 2144 10252 2208
rect 10316 2144 10332 2208
rect 10396 2144 10412 2208
rect 10476 2144 10492 2208
rect 10556 2144 10584 2208
rect 10224 274 10584 2144
rect 10224 38 10286 274
rect 10522 38 10584 274
rect 10224 -4 10584 38
rect 11524 14534 11884 15236
rect 14096 15194 14416 15236
rect 14096 14958 14138 15194
rect 14374 14958 14416 15194
rect 11524 14298 11586 14534
rect 11822 14298 11884 14534
rect 11524 12894 11884 14298
rect 11524 12658 11586 12894
rect 11822 12658 11884 12894
rect 11524 12544 11884 12658
rect 11524 12480 11552 12544
rect 11616 12480 11632 12544
rect 11696 12480 11712 12544
rect 11776 12480 11792 12544
rect 11856 12480 11884 12544
rect 11524 11456 11884 12480
rect 11524 11392 11552 11456
rect 11616 11392 11632 11456
rect 11696 11392 11712 11456
rect 11776 11392 11792 11456
rect 11856 11392 11884 11456
rect 11524 10894 11884 11392
rect 11524 10658 11586 10894
rect 11822 10658 11884 10894
rect 11524 10368 11884 10658
rect 11524 10304 11552 10368
rect 11616 10304 11632 10368
rect 11696 10304 11712 10368
rect 11776 10304 11792 10368
rect 11856 10304 11884 10368
rect 11524 9280 11884 10304
rect 11524 9216 11552 9280
rect 11616 9216 11632 9280
rect 11696 9216 11712 9280
rect 11776 9216 11792 9280
rect 11856 9216 11884 9280
rect 11524 8894 11884 9216
rect 11524 8658 11586 8894
rect 11822 8658 11884 8894
rect 11524 8192 11884 8658
rect 11524 8128 11552 8192
rect 11616 8128 11632 8192
rect 11696 8128 11712 8192
rect 11776 8128 11792 8192
rect 11856 8128 11884 8192
rect 11524 7104 11884 8128
rect 11524 7040 11552 7104
rect 11616 7040 11632 7104
rect 11696 7040 11712 7104
rect 11776 7040 11792 7104
rect 11856 7040 11884 7104
rect 11524 6894 11884 7040
rect 11524 6658 11586 6894
rect 11822 6658 11884 6894
rect 11524 6016 11884 6658
rect 11524 5952 11552 6016
rect 11616 5952 11632 6016
rect 11696 5952 11712 6016
rect 11776 5952 11792 6016
rect 11856 5952 11884 6016
rect 11524 4928 11884 5952
rect 11524 4864 11552 4928
rect 11616 4894 11632 4928
rect 11696 4894 11712 4928
rect 11776 4894 11792 4928
rect 11856 4864 11884 4928
rect 11524 4658 11586 4864
rect 11822 4658 11884 4864
rect 11524 3840 11884 4658
rect 11524 3776 11552 3840
rect 11616 3776 11632 3840
rect 11696 3776 11712 3840
rect 11776 3776 11792 3840
rect 11856 3776 11884 3840
rect 11524 2894 11884 3776
rect 11524 2752 11586 2894
rect 11822 2752 11884 2894
rect 11524 2688 11552 2752
rect 11856 2688 11884 2752
rect 11524 2658 11586 2688
rect 11822 2658 11884 2688
rect 11524 934 11884 2658
rect 11524 698 11586 934
rect 11822 698 11884 934
rect 11524 -4 11884 698
rect 13436 14534 13756 14576
rect 13436 14298 13478 14534
rect 13714 14298 13756 14534
rect 13436 12894 13756 14298
rect 13436 12658 13478 12894
rect 13714 12658 13756 12894
rect 13436 10894 13756 12658
rect 13436 10658 13478 10894
rect 13714 10658 13756 10894
rect 13436 8894 13756 10658
rect 13436 8658 13478 8894
rect 13714 8658 13756 8894
rect 13436 6894 13756 8658
rect 13436 6658 13478 6894
rect 13714 6658 13756 6894
rect 13436 4894 13756 6658
rect 13436 4658 13478 4894
rect 13714 4658 13756 4894
rect 13436 2894 13756 4658
rect 13436 2658 13478 2894
rect 13714 2658 13756 2894
rect 13436 934 13756 2658
rect 13436 698 13478 934
rect 13714 698 13756 934
rect 13436 656 13756 698
rect 14096 11594 14416 14958
rect 14096 11358 14138 11594
rect 14374 11358 14416 11594
rect 14096 9594 14416 11358
rect 14096 9358 14138 9594
rect 14374 9358 14416 9594
rect 14096 7594 14416 9358
rect 14096 7358 14138 7594
rect 14374 7358 14416 7594
rect 14096 5594 14416 7358
rect 14096 5358 14138 5594
rect 14374 5358 14416 5594
rect 14096 3594 14416 5358
rect 14096 3358 14138 3594
rect 14374 3358 14416 3594
rect 14096 274 14416 3358
rect 14096 38 14138 274
rect 14374 38 14416 274
rect 14096 -4 14416 38
<< via4 >>
rect -1034 14958 -798 15194
rect -1034 11358 -798 11594
rect -1034 9358 -798 9594
rect -1034 7358 -798 7594
rect -1034 5358 -798 5594
rect -1034 3358 -798 3594
rect -374 14298 -138 14534
rect -374 12658 -138 12894
rect -374 10658 -138 10894
rect -374 8658 -138 8894
rect -374 6658 -138 6894
rect -374 4658 -138 4894
rect -374 2658 -138 2894
rect -374 698 -138 934
rect 1586 14298 1822 14534
rect 1586 12658 1822 12894
rect 1586 10658 1822 10894
rect 1586 8658 1822 8894
rect 1586 6658 1822 6894
rect 1586 4864 1616 4894
rect 1616 4864 1632 4894
rect 1632 4864 1696 4894
rect 1696 4864 1712 4894
rect 1712 4864 1776 4894
rect 1776 4864 1792 4894
rect 1792 4864 1822 4894
rect 1586 4658 1822 4864
rect 1586 2752 1822 2894
rect 1586 2688 1616 2752
rect 1616 2688 1632 2752
rect 1632 2688 1696 2752
rect 1696 2688 1712 2752
rect 1712 2688 1776 2752
rect 1776 2688 1792 2752
rect 1792 2688 1822 2752
rect 1586 2658 1822 2688
rect 1586 698 1822 934
rect -1034 38 -798 274
rect 2286 14958 2522 15194
rect 2286 11358 2522 11594
rect 2286 9358 2522 9594
rect 2286 7584 2316 7594
rect 2316 7584 2332 7594
rect 2332 7584 2396 7594
rect 2396 7584 2412 7594
rect 2412 7584 2476 7594
rect 2476 7584 2492 7594
rect 2492 7584 2522 7594
rect 2286 7358 2522 7584
rect 2286 5472 2522 5594
rect 2286 5408 2316 5472
rect 2316 5408 2332 5472
rect 2332 5408 2396 5472
rect 2396 5408 2412 5472
rect 2412 5408 2476 5472
rect 2476 5408 2492 5472
rect 2492 5408 2522 5472
rect 2286 5358 2522 5408
rect 2286 3358 2522 3594
rect 2286 38 2522 274
rect 3586 14298 3822 14534
rect 3586 12658 3822 12894
rect 3586 10658 3822 10894
rect 3586 8658 3822 8894
rect 3586 6658 3822 6894
rect 3586 4864 3616 4894
rect 3616 4864 3632 4894
rect 3632 4864 3696 4894
rect 3696 4864 3712 4894
rect 3712 4864 3776 4894
rect 3776 4864 3792 4894
rect 3792 4864 3822 4894
rect 3586 4658 3822 4864
rect 3586 2752 3822 2894
rect 3586 2688 3616 2752
rect 3616 2688 3632 2752
rect 3632 2688 3696 2752
rect 3696 2688 3712 2752
rect 3712 2688 3776 2752
rect 3776 2688 3792 2752
rect 3792 2688 3822 2752
rect 3586 2658 3822 2688
rect 3586 698 3822 934
rect 4286 14958 4522 15194
rect 4286 11358 4522 11594
rect 4286 9358 4522 9594
rect 4286 7584 4316 7594
rect 4316 7584 4332 7594
rect 4332 7584 4396 7594
rect 4396 7584 4412 7594
rect 4412 7584 4476 7594
rect 4476 7584 4492 7594
rect 4492 7584 4522 7594
rect 4286 7358 4522 7584
rect 4286 5472 4522 5594
rect 4286 5408 4316 5472
rect 4316 5408 4332 5472
rect 4332 5408 4396 5472
rect 4396 5408 4412 5472
rect 4412 5408 4476 5472
rect 4476 5408 4492 5472
rect 4492 5408 4522 5472
rect 4286 5358 4522 5408
rect 4286 3358 4522 3594
rect 4286 38 4522 274
rect 5586 14298 5822 14534
rect 5586 12658 5822 12894
rect 5586 10658 5822 10894
rect 5586 8658 5822 8894
rect 5586 6658 5822 6894
rect 5586 4864 5616 4894
rect 5616 4864 5632 4894
rect 5632 4864 5696 4894
rect 5696 4864 5712 4894
rect 5712 4864 5776 4894
rect 5776 4864 5792 4894
rect 5792 4864 5822 4894
rect 5586 4658 5822 4864
rect 5586 2752 5822 2894
rect 5586 2688 5616 2752
rect 5616 2688 5632 2752
rect 5632 2688 5696 2752
rect 5696 2688 5712 2752
rect 5712 2688 5776 2752
rect 5776 2688 5792 2752
rect 5792 2688 5822 2752
rect 5586 2658 5822 2688
rect 5586 698 5822 934
rect 6286 14958 6522 15194
rect 6286 11358 6522 11594
rect 6286 9358 6522 9594
rect 6286 7584 6316 7594
rect 6316 7584 6332 7594
rect 6332 7584 6396 7594
rect 6396 7584 6412 7594
rect 6412 7584 6476 7594
rect 6476 7584 6492 7594
rect 6492 7584 6522 7594
rect 6286 7358 6522 7584
rect 6286 5472 6522 5594
rect 6286 5408 6316 5472
rect 6316 5408 6332 5472
rect 6332 5408 6396 5472
rect 6396 5408 6412 5472
rect 6412 5408 6476 5472
rect 6476 5408 6492 5472
rect 6492 5408 6522 5472
rect 6286 5358 6522 5408
rect 6286 3358 6522 3594
rect 6286 38 6522 274
rect 7586 14298 7822 14534
rect 7586 12658 7822 12894
rect 7586 10658 7822 10894
rect 7586 8658 7822 8894
rect 7586 6658 7822 6894
rect 7586 4864 7616 4894
rect 7616 4864 7632 4894
rect 7632 4864 7696 4894
rect 7696 4864 7712 4894
rect 7712 4864 7776 4894
rect 7776 4864 7792 4894
rect 7792 4864 7822 4894
rect 7586 4658 7822 4864
rect 7586 2752 7822 2894
rect 7586 2688 7616 2752
rect 7616 2688 7632 2752
rect 7632 2688 7696 2752
rect 7696 2688 7712 2752
rect 7712 2688 7776 2752
rect 7776 2688 7792 2752
rect 7792 2688 7822 2752
rect 7586 2658 7822 2688
rect 7586 698 7822 934
rect 8286 14958 8522 15194
rect 8286 11358 8522 11594
rect 8286 9358 8522 9594
rect 8286 7584 8316 7594
rect 8316 7584 8332 7594
rect 8332 7584 8396 7594
rect 8396 7584 8412 7594
rect 8412 7584 8476 7594
rect 8476 7584 8492 7594
rect 8492 7584 8522 7594
rect 8286 7358 8522 7584
rect 8286 5472 8522 5594
rect 8286 5408 8316 5472
rect 8316 5408 8332 5472
rect 8332 5408 8396 5472
rect 8396 5408 8412 5472
rect 8412 5408 8476 5472
rect 8476 5408 8492 5472
rect 8492 5408 8522 5472
rect 8286 5358 8522 5408
rect 8286 3358 8522 3594
rect 8286 38 8522 274
rect 9586 14298 9822 14534
rect 9586 12658 9822 12894
rect 9586 10658 9822 10894
rect 9586 8658 9822 8894
rect 9586 6658 9822 6894
rect 9586 4864 9616 4894
rect 9616 4864 9632 4894
rect 9632 4864 9696 4894
rect 9696 4864 9712 4894
rect 9712 4864 9776 4894
rect 9776 4864 9792 4894
rect 9792 4864 9822 4894
rect 9586 4658 9822 4864
rect 9586 2752 9822 2894
rect 9586 2688 9616 2752
rect 9616 2688 9632 2752
rect 9632 2688 9696 2752
rect 9696 2688 9712 2752
rect 9712 2688 9776 2752
rect 9776 2688 9792 2752
rect 9792 2688 9822 2752
rect 9586 2658 9822 2688
rect 9586 698 9822 934
rect 10286 14958 10522 15194
rect 10286 11358 10522 11594
rect 10286 9358 10522 9594
rect 10286 7584 10316 7594
rect 10316 7584 10332 7594
rect 10332 7584 10396 7594
rect 10396 7584 10412 7594
rect 10412 7584 10476 7594
rect 10476 7584 10492 7594
rect 10492 7584 10522 7594
rect 10286 7358 10522 7584
rect 10286 5472 10522 5594
rect 10286 5408 10316 5472
rect 10316 5408 10332 5472
rect 10332 5408 10396 5472
rect 10396 5408 10412 5472
rect 10412 5408 10476 5472
rect 10476 5408 10492 5472
rect 10492 5408 10522 5472
rect 10286 5358 10522 5408
rect 10286 3358 10522 3594
rect 10286 38 10522 274
rect 14138 14958 14374 15194
rect 11586 14298 11822 14534
rect 11586 12658 11822 12894
rect 11586 10658 11822 10894
rect 11586 8658 11822 8894
rect 11586 6658 11822 6894
rect 11586 4864 11616 4894
rect 11616 4864 11632 4894
rect 11632 4864 11696 4894
rect 11696 4864 11712 4894
rect 11712 4864 11776 4894
rect 11776 4864 11792 4894
rect 11792 4864 11822 4894
rect 11586 4658 11822 4864
rect 11586 2752 11822 2894
rect 11586 2688 11616 2752
rect 11616 2688 11632 2752
rect 11632 2688 11696 2752
rect 11696 2688 11712 2752
rect 11712 2688 11776 2752
rect 11776 2688 11792 2752
rect 11792 2688 11822 2752
rect 11586 2658 11822 2688
rect 11586 698 11822 934
rect 13478 14298 13714 14534
rect 13478 12658 13714 12894
rect 13478 10658 13714 10894
rect 13478 8658 13714 8894
rect 13478 6658 13714 6894
rect 13478 4658 13714 4894
rect 13478 2658 13714 2894
rect 13478 698 13714 934
rect 14138 11358 14374 11594
rect 14138 9358 14374 9594
rect 14138 7358 14374 7594
rect 14138 5358 14374 5594
rect 14138 3358 14374 3594
rect 14138 38 14374 274
<< metal5 >>
rect -1076 15194 14416 15236
rect -1076 14958 -1034 15194
rect -798 14958 2286 15194
rect 2522 14958 4286 15194
rect 4522 14958 6286 15194
rect 6522 14958 8286 15194
rect 8522 14958 10286 15194
rect 10522 14958 14138 15194
rect 14374 14958 14416 15194
rect -1076 14916 14416 14958
rect -416 14534 13756 14576
rect -416 14298 -374 14534
rect -138 14298 1586 14534
rect 1822 14298 3586 14534
rect 3822 14298 5586 14534
rect 5822 14298 7586 14534
rect 7822 14298 9586 14534
rect 9822 14298 11586 14534
rect 11822 14298 13478 14534
rect 13714 14298 13756 14534
rect -416 14256 13756 14298
rect -1076 12894 14416 12956
rect -1076 12658 -374 12894
rect -138 12658 1586 12894
rect 1822 12658 3586 12894
rect 3822 12658 5586 12894
rect 5822 12658 7586 12894
rect 7822 12658 9586 12894
rect 9822 12658 11586 12894
rect 11822 12658 13478 12894
rect 13714 12658 14416 12894
rect -1076 12596 14416 12658
rect -1076 11594 14416 11656
rect -1076 11358 -1034 11594
rect -798 11358 2286 11594
rect 2522 11358 4286 11594
rect 4522 11358 6286 11594
rect 6522 11358 8286 11594
rect 8522 11358 10286 11594
rect 10522 11358 14138 11594
rect 14374 11358 14416 11594
rect -1076 11296 14416 11358
rect -1076 10894 14416 10956
rect -1076 10658 -374 10894
rect -138 10658 1586 10894
rect 1822 10658 3586 10894
rect 3822 10658 5586 10894
rect 5822 10658 7586 10894
rect 7822 10658 9586 10894
rect 9822 10658 11586 10894
rect 11822 10658 13478 10894
rect 13714 10658 14416 10894
rect -1076 10596 14416 10658
rect -1076 9594 14416 9656
rect -1076 9358 -1034 9594
rect -798 9358 2286 9594
rect 2522 9358 4286 9594
rect 4522 9358 6286 9594
rect 6522 9358 8286 9594
rect 8522 9358 10286 9594
rect 10522 9358 14138 9594
rect 14374 9358 14416 9594
rect -1076 9296 14416 9358
rect -1076 8894 14416 8956
rect -1076 8658 -374 8894
rect -138 8658 1586 8894
rect 1822 8658 3586 8894
rect 3822 8658 5586 8894
rect 5822 8658 7586 8894
rect 7822 8658 9586 8894
rect 9822 8658 11586 8894
rect 11822 8658 13478 8894
rect 13714 8658 14416 8894
rect -1076 8596 14416 8658
rect -1076 7594 14416 7656
rect -1076 7358 -1034 7594
rect -798 7358 2286 7594
rect 2522 7358 4286 7594
rect 4522 7358 6286 7594
rect 6522 7358 8286 7594
rect 8522 7358 10286 7594
rect 10522 7358 14138 7594
rect 14374 7358 14416 7594
rect -1076 7296 14416 7358
rect -1076 6894 14416 6956
rect -1076 6658 -374 6894
rect -138 6658 1586 6894
rect 1822 6658 3586 6894
rect 3822 6658 5586 6894
rect 5822 6658 7586 6894
rect 7822 6658 9586 6894
rect 9822 6658 11586 6894
rect 11822 6658 13478 6894
rect 13714 6658 14416 6894
rect -1076 6596 14416 6658
rect -1076 5594 14416 5656
rect -1076 5358 -1034 5594
rect -798 5358 2286 5594
rect 2522 5358 4286 5594
rect 4522 5358 6286 5594
rect 6522 5358 8286 5594
rect 8522 5358 10286 5594
rect 10522 5358 14138 5594
rect 14374 5358 14416 5594
rect -1076 5296 14416 5358
rect -1076 4894 14416 4956
rect -1076 4658 -374 4894
rect -138 4658 1586 4894
rect 1822 4658 3586 4894
rect 3822 4658 5586 4894
rect 5822 4658 7586 4894
rect 7822 4658 9586 4894
rect 9822 4658 11586 4894
rect 11822 4658 13478 4894
rect 13714 4658 14416 4894
rect -1076 4596 14416 4658
rect -1076 3594 14416 3656
rect -1076 3358 -1034 3594
rect -798 3358 2286 3594
rect 2522 3358 4286 3594
rect 4522 3358 6286 3594
rect 6522 3358 8286 3594
rect 8522 3358 10286 3594
rect 10522 3358 14138 3594
rect 14374 3358 14416 3594
rect -1076 3296 14416 3358
rect -1076 2894 14416 2956
rect -1076 2658 -374 2894
rect -138 2658 1586 2894
rect 1822 2658 3586 2894
rect 3822 2658 5586 2894
rect 5822 2658 7586 2894
rect 7822 2658 9586 2894
rect 9822 2658 11586 2894
rect 11822 2658 13478 2894
rect 13714 2658 14416 2894
rect -1076 2596 14416 2658
rect -416 934 13756 976
rect -416 698 -374 934
rect -138 698 1586 934
rect 1822 698 3586 934
rect 3822 698 5586 934
rect 5822 698 7586 934
rect 7822 698 9586 934
rect 9822 698 11586 934
rect 11822 698 13478 934
rect 13714 698 13756 934
rect -416 656 13756 698
rect -1076 274 14416 316
rect -1076 38 -1034 274
rect -798 38 2286 274
rect 2522 38 4286 274
rect 4522 38 6286 274
rect 6522 38 8286 274
rect 8522 38 10286 274
rect 10522 38 14138 274
rect 14374 38 14416 274
rect -1076 -4 14416 38
use sky130_fd_sc_hd__inv_2  _066_
timestamp -28799
transform -1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _067_
timestamp -28799
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _068_
timestamp -28799
transform 1 0 5336 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _069_
timestamp -28799
transform 1 0 6624 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _070_
timestamp -28799
transform 1 0 5704 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _071_
timestamp -28799
transform 1 0 5152 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _072_
timestamp -28799
transform -1 0 5704 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _073_
timestamp -28799
transform 1 0 4600 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _074_
timestamp -28799
transform 1 0 3956 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _075_
timestamp -28799
transform -1 0 2116 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _076_
timestamp -28799
transform -1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _077_
timestamp -28799
transform 1 0 5520 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _078_
timestamp -28799
transform -1 0 4232 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _079_
timestamp -28799
transform 1 0 3036 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _080_
timestamp -28799
transform 1 0 2300 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _081_
timestamp -28799
transform -1 0 3680 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _082_
timestamp -28799
transform 1 0 1840 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _083_
timestamp -28799
transform -1 0 2300 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _084_
timestamp -28799
transform 1 0 1472 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _085_
timestamp -28799
transform 1 0 1932 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _086_
timestamp -28799
transform 1 0 3036 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _087_
timestamp -28799
transform 1 0 2668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _088_
timestamp -28799
transform -1 0 4232 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _089_
timestamp -28799
transform -1 0 2576 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _090_
timestamp -28799
transform 1 0 3680 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _091_
timestamp -28799
transform 1 0 4876 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _092_
timestamp -28799
transform 1 0 2116 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _093_
timestamp -28799
transform -1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _094_
timestamp -28799
transform -1 0 5520 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _095_
timestamp -28799
transform -1 0 8280 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _096_
timestamp -28799
transform 1 0 5520 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _097_
timestamp -28799
transform 1 0 6348 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _098_
timestamp -28799
transform 1 0 6072 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _099_
timestamp -28799
transform -1 0 6256 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _100_
timestamp -28799
transform 1 0 5244 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _101_
timestamp -28799
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _102_
timestamp -28799
transform -1 0 7728 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _103_
timestamp -28799
transform -1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _104_
timestamp -28799
transform -1 0 10212 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _105_
timestamp -28799
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _106_
timestamp -28799
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _107_
timestamp -28799
transform -1 0 8740 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _108_
timestamp -28799
transform 1 0 7820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _109_
timestamp -28799
transform -1 0 11408 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _110_
timestamp -28799
transform 1 0 9660 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _111_
timestamp -28799
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _112_
timestamp -28799
transform -1 0 9568 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _113_
timestamp -28799
transform -1 0 11408 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _114_
timestamp -28799
transform -1 0 10304 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _115_
timestamp -28799
transform 1 0 10028 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _116_
timestamp -28799
transform 1 0 11500 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _117_
timestamp -28799
transform 1 0 10304 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _118_
timestamp -28799
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _119_
timestamp -28799
transform -1 0 10948 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _120_
timestamp -28799
transform 1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _121_
timestamp -28799
transform -1 0 9568 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _122_
timestamp -28799
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _123_
timestamp -28799
transform -1 0 11040 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _124_
timestamp -28799
transform -1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _125_
timestamp -28799
transform -1 0 11960 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _126_
timestamp -28799
transform -1 0 10580 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _127_
timestamp -28799
transform -1 0 9200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _128_
timestamp -28799
transform -1 0 11224 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _129_
timestamp -28799
transform -1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _130_
timestamp -28799
transform -1 0 9844 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _131_
timestamp -28799
transform 1 0 9016 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _132_
timestamp -28799
transform -1 0 8832 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _133_
timestamp -28799
transform -1 0 7360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _134_
timestamp -28799
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp -28799
transform 1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp -28799
transform -1 0 3588 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp -28799
transform -1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp -28799
transform -1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp -28799
transform -1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp -28799
transform -1 0 3956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp -28799
transform 1 0 3956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp -28799
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp -28799
transform -1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp -28799
transform -1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp -28799
transform -1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp -28799
transform -1 0 8648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp -28799
transform -1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp -28799
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp -28799
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _150_
timestamp -28799
transform 1 0 7636 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp -28799
transform -1 0 9568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152_
timestamp -28799
transform 1 0 9384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _153_
timestamp -28799
transform 1 0 9752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp -28799
transform -1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp -28799
transform 1 0 10672 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp -28799
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp -28799
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp -28799
transform 1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp -28799
transform -1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp -28799
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp -28799
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _162_
timestamp -28799
transform 1 0 3036 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _163_
timestamp -28799
transform -1 0 7084 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _164_
timestamp -28799
transform -1 0 8188 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _165_
timestamp -28799
transform 1 0 3864 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _166_
timestamp -28799
transform 1 0 1472 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _167_
timestamp -28799
transform -1 0 3680 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _168_
timestamp -28799
transform 1 0 3772 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _169_
timestamp -28799
transform 1 0 1472 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _170_
timestamp -28799
transform 1 0 1840 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _171_
timestamp -28799
transform -1 0 5612 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _172_
timestamp -28799
transform 1 0 1840 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _173_
timestamp -28799
transform 1 0 2852 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _174_
timestamp -28799
transform 1 0 4140 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _175_
timestamp -28799
transform 1 0 5980 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _176_
timestamp -28799
transform 1 0 6716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _177_
timestamp -28799
transform 1 0 5612 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _178_
timestamp -28799
transform 1 0 6992 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _179_
timestamp -28799
transform 1 0 6992 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _180_
timestamp -28799
transform 1 0 6992 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _181_
timestamp -28799
transform 1 0 7912 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _182_
timestamp -28799
transform 1 0 8464 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _183_
timestamp -28799
transform 1 0 10120 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _184_
timestamp -28799
transform 1 0 9568 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _185_
timestamp -28799
transform 1 0 10120 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _186_
timestamp -28799
transform 1 0 7912 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _187_
timestamp -28799
transform 1 0 9936 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _188_
timestamp -28799
transform 1 0 9568 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _189_
timestamp -28799
transform 1 0 9660 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _190_
timestamp -28799
transform 1 0 9568 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _191_
timestamp -28799
transform 1 0 7636 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -28799
transform 1 0 5152 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp -28799
transform -1 0 6072 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp -28799
transform 1 0 8924 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp -28799
transform -1 0 5612 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp -28799
transform 1 0 8924 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp -28799
transform 1 0 4232 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload1
timestamp -28799
transform 1 0 8924 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload2
timestamp -28799
transform 1 0 3772 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout32
timestamp -28799
transform -1 0 8648 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp -28799
transform -1 0 11408 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout34
timestamp -28799
transform 1 0 9200 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp -28799
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636939656
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15
timestamp -28799
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp -28799
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp -28799
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38
timestamp 1636939656
transform 1 0 4600 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50
timestamp -28799
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp -28799
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88
timestamp -28799
transform 1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp -28799
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp -28799
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp -28799
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_16
timestamp -28799
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp -28799
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -28799
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_70
timestamp -28799
transform 1 0 7544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_91
timestamp -28799
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_116
timestamp -28799
transform 1 0 11776 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp -28799
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp -28799
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp -28799
transform 1 0 4048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_78
timestamp -28799
transform 1 0 8280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp -28799
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp -28799
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_113
timestamp -28799
transform 1 0 11500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp -28799
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_45
timestamp -28799
transform 1 0 5244 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_65
timestamp -28799
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp -28799
transform 1 0 8648 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -28799
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp -28799
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636939656
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_15
timestamp -28799
transform 1 0 2484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp -28799
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp -28799
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_11
timestamp -28799
transform 1 0 2116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_25
timestamp -28799
transform 1 0 3404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_35
timestamp -28799
transform 1 0 4324 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp -28799
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp -28799
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_65
timestamp -28799
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_73
timestamp -28799
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp -28799
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp -28799
transform 1 0 8464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_103
timestamp -28799
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp -28799
transform 1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_14
timestamp -28799
transform 1 0 2392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_34
timestamp -28799
transform 1 0 4232 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_40
timestamp -28799
transform 1 0 4784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp -28799
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp -28799
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636939656
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636939656
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_81
timestamp -28799
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp -28799
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp -28799
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_13
timestamp 1636939656
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp -28799
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636939656
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636939656
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636939656
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_72
timestamp 1636939656
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_92
timestamp -28799
transform 1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp -28799
transform 1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp -28799
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636939656
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636939656
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp -28799
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -28799
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_57
timestamp -28799
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_63
timestamp -28799
transform 1 0 6900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_95
timestamp -28799
transform 1 0 9844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_117
timestamp -28799
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_7
timestamp -28799
transform 1 0 1748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp -28799
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636939656
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp -28799
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp -28799
transform 1 0 9200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_96
timestamp -28799
transform 1 0 9936 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp -28799
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_16
timestamp -28799
transform 1 0 2576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_20
timestamp -28799
transform 1 0 2944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_28
timestamp -28799
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp -28799
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636939656
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_69
timestamp -28799
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_77
timestamp -28799
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_107
timestamp -28799
transform 1 0 10948 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp -28799
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp -28799
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_61
timestamp -28799
transform 1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp -28799
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_25
timestamp -28799
transform 1 0 3404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp -28799
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp -28799
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636939656
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_69
timestamp -28799
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_102
timestamp -28799
transform 1 0 10488 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp -28799
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp -28799
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp -28799
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp -28799
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp -28799
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_34
timestamp -28799
transform 1 0 4232 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_43
timestamp 1636939656
transform 1 0 5060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_55
timestamp 1636939656
transform 1 0 6164 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_67
timestamp -28799
transform 1 0 7268 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp -28799
transform 1 0 11776 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_7
timestamp 1636939656
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_19
timestamp -28799
transform 1 0 2852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp -28799
transform 1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp -28799
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636939656
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp -28799
transform 1 0 7452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_77
timestamp -28799
transform 1 0 8188 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_83
timestamp -28799
transform 1 0 8740 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636939656
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636939656
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp -28799
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp -28799
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp -28799
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_68
timestamp 1636939656
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp -28799
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_92
timestamp -28799
transform 1 0 9568 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636939656
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp -28799
transform 1 0 2484 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_41
timestamp -28799
transform 1 0 4876 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp -28799
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_77
timestamp -28799
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp -28799
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636939656
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636939656
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -28799
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp -28799
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_37
timestamp -28799
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_49
timestamp -28799
transform 1 0 5612 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_68
timestamp 1636939656
transform 1 0 7360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp -28799
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp -28799
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp -28799
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp -28799
transform 1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_108
timestamp -28799
transform 1 0 11040 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp -28799
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636939656
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636939656
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_27
timestamp -28799
transform 1 0 3588 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_29
timestamp -28799
transform 1 0 3772 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_35
timestamp -28799
transform 1 0 4324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_51
timestamp -28799
transform 1 0 5796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp -28799
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_63
timestamp 1636939656
transform 1 0 6900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_75
timestamp -28799
transform 1 0 8004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_83
timestamp -28799
transform 1 0 8740 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_85
timestamp -28799
transform 1 0 8924 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp -28799
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -28799
transform -1 0 10120 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -28799
transform -1 0 11592 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -28799
transform -1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp -28799
transform -1 0 5336 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp -28799
transform -1 0 4232 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp -28799
transform -1 0 3496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp -28799
transform -1 0 7544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp -28799
transform -1 0 8096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp -28799
transform -1 0 5520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp -28799
transform -1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp -28799
transform -1 0 3312 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp -28799
transform -1 0 6624 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp -28799
transform -1 0 3404 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp -28799
transform -1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp -28799
transform -1 0 8188 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp -28799
transform -1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp -28799
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp -28799
transform -1 0 11040 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp -28799
transform -1 0 9568 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp -28799
transform -1 0 9568 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp -28799
transform -1 0 9200 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp -28799
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp -28799
transform -1 0 11316 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp -28799
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp -28799
transform -1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp -28799
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  MIPSpipeline_36
timestamp -28799
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  MIPSpipeline_37
timestamp -28799
transform 1 0 9476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -28799
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -28799
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -28799
transform -1 0 3680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -28799
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -28799
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -28799
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -28799
transform -1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -28799
transform -1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -28799
transform 1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -28799
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -28799
transform 1 0 11592 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -28799
transform 1 0 11592 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -28799
transform 1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -28799
transform 1 0 11592 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -28799
transform 1 0 11408 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -28799
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -28799
transform 1 0 11592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -28799
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -28799
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -28799
transform 1 0 11592 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -28799
transform -1 0 4784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -28799
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -28799
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -28799
transform 1 0 4784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -28799
transform 1 0 6532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -28799
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -28799
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -28799
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -28799
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -28799
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_20
timestamp -28799
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -28799
transform -1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_21
timestamp -28799
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -28799
transform -1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_22
timestamp -28799
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -28799
transform -1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_23
timestamp -28799
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -28799
transform -1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_24
timestamp -28799
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -28799
transform -1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_25
timestamp -28799
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -28799
transform -1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_26
timestamp -28799
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -28799
transform -1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_27
timestamp -28799
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -28799
transform -1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_28
timestamp -28799
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -28799
transform -1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_29
timestamp -28799
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -28799
transform -1 0 12236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_30
timestamp -28799
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -28799
transform -1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_31
timestamp -28799
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -28799
transform -1 0 12236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_32
timestamp -28799
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -28799
transform -1 0 12236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_33
timestamp -28799
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -28799
transform -1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_34
timestamp -28799
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -28799
transform -1 0 12236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_35
timestamp -28799
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -28799
transform -1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_36
timestamp -28799
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -28799
transform -1 0 12236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_37
timestamp -28799
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -28799
transform -1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_38
timestamp -28799
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -28799
transform -1 0 12236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_39
timestamp -28799
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -28799
transform -1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_40
timestamp -28799
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_41
timestamp -28799
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_42
timestamp -28799
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_43
timestamp -28799
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -28799
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp -28799
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -28799
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -28799
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_48
timestamp -28799
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_49
timestamp -28799
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_50
timestamp -28799
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_51
timestamp -28799
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_52
timestamp -28799
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_53
timestamp -28799
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_54
timestamp -28799
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_55
timestamp -28799
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_56
timestamp -28799
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_57
timestamp -28799
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_58
timestamp -28799
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_59
timestamp -28799
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_60
timestamp -28799
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_61
timestamp -28799
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_62
timestamp -28799
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_63
timestamp -28799
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_64
timestamp -28799
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_65
timestamp -28799
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_66
timestamp -28799
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_67
timestamp -28799
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_68
timestamp -28799
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_69
timestamp -28799
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_70
timestamp -28799
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_71
timestamp -28799
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_72
timestamp -28799
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_73
timestamp -28799
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_74
timestamp -28799
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_75
timestamp -28799
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_76
timestamp -28799
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_77
timestamp -28799
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_78
timestamp -28799
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_79
timestamp -28799
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_80
timestamp -28799
transform 1 0 3680 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_81
timestamp -28799
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_82
timestamp -28799
transform 1 0 8832 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_83
timestamp -28799
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
<< labels >>
flabel metal4 s -1076 -4 -756 15236 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -1076 -4 14416 316 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -1076 14916 14416 15236 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14096 -4 14416 15236 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2224 -4 2584 15236 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4224 -4 4584 15236 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6224 -4 6584 15236 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8224 -4 8584 15236 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10224 -4 10584 15236 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -1076 3296 14416 3656 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -1076 5296 14416 5656 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -1076 7296 14416 7656 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -1076 9296 14416 9656 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -1076 11296 14416 11656 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s -416 656 -96 14576 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -416 656 13756 976 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -416 14256 13756 14576 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13436 656 13756 14576 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 1524 -4 1884 15236 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3524 -4 3884 15236 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5524 -4 5884 15236 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7524 -4 7884 15236 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9524 -4 9884 15236 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11524 -4 11884 15236 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -1076 2596 14416 2956 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -1076 4596 14416 4956 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -1076 6596 14416 6956 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -1076 8596 14416 8956 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -1076 10596 14416 10956 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -1076 12596 14416 12956 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 12607 2728 13407 2848 0 FreeSans 480 0 0 0 current_pc[0]
port 3 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 current_pc[10]
port 4 nsew signal output
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 current_pc[11]
port 5 nsew signal output
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 current_pc[12]
port 6 nsew signal output
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 current_pc[13]
port 7 nsew signal output
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 current_pc[14]
port 8 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 current_pc[15]
port 9 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 current_pc[16]
port 10 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 current_pc[17]
port 11 nsew signal output
flabel metal3 s 12607 7488 13407 7608 0 FreeSans 480 0 0 0 current_pc[18]
port 12 nsew signal output
flabel metal3 s 12607 8168 13407 8288 0 FreeSans 480 0 0 0 current_pc[19]
port 13 nsew signal output
flabel metal3 s 12607 12928 13407 13048 0 FreeSans 480 0 0 0 current_pc[1]
port 14 nsew signal output
flabel metal3 s 12607 9528 13407 9648 0 FreeSans 480 0 0 0 current_pc[20]
port 15 nsew signal output
flabel metal3 s 12607 10888 13407 11008 0 FreeSans 480 0 0 0 current_pc[21]
port 16 nsew signal output
flabel metal3 s 12607 12248 13407 12368 0 FreeSans 480 0 0 0 current_pc[22]
port 17 nsew signal output
flabel metal3 s 12607 11568 13407 11688 0 FreeSans 480 0 0 0 current_pc[23]
port 18 nsew signal output
flabel metal3 s 12607 10208 13407 10328 0 FreeSans 480 0 0 0 current_pc[24]
port 19 nsew signal output
flabel metal3 s 12607 8848 13407 8968 0 FreeSans 480 0 0 0 current_pc[25]
port 20 nsew signal output
flabel metal3 s 12607 6128 13407 6248 0 FreeSans 480 0 0 0 current_pc[26]
port 21 nsew signal output
flabel metal3 s 12607 6808 13407 6928 0 FreeSans 480 0 0 0 current_pc[27]
port 22 nsew signal output
flabel metal3 s 12607 5448 13407 5568 0 FreeSans 480 0 0 0 current_pc[28]
port 23 nsew signal output
flabel metal3 s 12607 4088 13407 4208 0 FreeSans 480 0 0 0 current_pc[29]
port 24 nsew signal output
flabel metal2 s 4526 14751 4582 15551 0 FreeSans 224 90 0 0 current_pc[2]
port 25 nsew signal output
flabel metal3 s 12607 3408 13407 3528 0 FreeSans 480 0 0 0 current_pc[30]
port 26 nsew signal output
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 current_pc[31]
port 27 nsew signal output
flabel metal2 s 5170 14751 5226 15551 0 FreeSans 224 90 0 0 current_pc[3]
port 28 nsew signal output
flabel metal2 s 6458 14751 6514 15551 0 FreeSans 224 90 0 0 current_pc[4]
port 29 nsew signal output
flabel metal2 s 5814 14751 5870 15551 0 FreeSans 224 90 0 0 current_pc[5]
port 30 nsew signal output
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 current_pc[6]
port 31 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 current_pc[7]
port 32 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 current_pc[8]
port 33 nsew signal output
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 current_pc[9]
port 34 nsew signal output
flabel metal3 s 12607 4768 13407 4888 0 FreeSans 480 0 0 0 reset
port 35 nsew signal input
rlabel metal1 6670 13056 6670 13056 0 VGND
rlabel metal1 6670 12512 6670 12512 0 VPWR
rlabel metal1 2116 5134 2116 5134 0 PC4\[10\]
rlabel metal1 4232 5746 4232 5746 0 PC4\[11\]
rlabel metal1 2070 2958 2070 2958 0 PC4\[12\]
rlabel metal2 2714 3536 2714 3536 0 PC4\[13\]
rlabel metal1 4830 2958 4830 2958 0 PC4\[14\]
rlabel metal1 6072 2822 6072 2822 0 PC4\[15\]
rlabel metal1 6900 4522 6900 4522 0 PC4\[16\]
rlabel metal1 6164 5338 6164 5338 0 PC4\[17\]
rlabel metal1 7222 6970 7222 6970 0 PC4\[18\]
rlabel metal2 7314 8092 7314 8092 0 PC4\[19\]
rlabel metal2 7314 9452 7314 9452 0 PC4\[20\]
rlabel metal2 8234 9588 8234 9588 0 PC4\[21\]
rlabel metal1 8878 11322 8878 11322 0 PC4\[22\]
rlabel metal1 10120 12614 10120 12614 0 PC4\[23\]
rlabel metal1 10258 10574 10258 10574 0 PC4\[24\]
rlabel metal1 9706 8058 9706 8058 0 PC4\[25\]
rlabel metal2 8970 5984 8970 5984 0 PC4\[26\]
rlabel metal1 10028 5338 10028 5338 0 PC4\[27\]
rlabel metal1 10028 5882 10028 5882 0 PC4\[28\]
rlabel metal1 10028 3434 10028 3434 0 PC4\[29\]
rlabel metal1 3358 11832 3358 11832 0 PC4\[2\]
rlabel metal2 9890 3196 9890 3196 0 PC4\[30\]
rlabel metal1 8096 2618 8096 2618 0 PC4\[31\]
rlabel metal1 6440 11186 6440 11186 0 PC4\[3\]
rlabel metal1 6578 12682 6578 12682 0 PC4\[4\]
rlabel metal1 4416 10574 4416 10574 0 PC4\[5\]
rlabel metal1 1656 9622 1656 9622 0 PC4\[6\]
rlabel metal2 3358 9418 3358 9418 0 PC4\[7\]
rlabel metal1 3634 8364 3634 8364 0 PC4\[8\]
rlabel metal1 1886 6970 1886 6970 0 PC4\[9\]
rlabel metal2 4094 11934 4094 11934 0 _000_
rlabel metal1 6493 11050 6493 11050 0 _001_
rlabel metal2 7222 11934 7222 11934 0 _002_
rlabel metal2 4922 10472 4922 10472 0 _003_
rlabel metal1 3227 9622 3227 9622 0 _004_
rlabel metal2 2898 9010 2898 9010 0 _005_
rlabel metal1 5527 8534 5527 8534 0 _006_
rlabel metal1 3227 7446 3227 7446 0 _007_
rlabel metal1 3634 6086 3634 6086 0 _008_
rlabel metal1 4140 6086 4140 6086 0 _009_
rlabel metal1 3641 3434 3641 3434 0 _010_
rlabel metal1 4423 3094 4423 3094 0 _011_
rlabel metal2 5198 3672 5198 3672 0 _012_
rlabel metal1 7544 2618 7544 2618 0 _013_
rlabel metal1 8326 3706 8326 3706 0 _014_
rlabel metal1 7367 5610 7367 5610 0 _015_
rlabel metal1 9115 7446 9115 7446 0 _016_
rlabel metal1 9161 7786 9161 7786 0 _017_
rlabel metal1 7866 9350 7866 9350 0 _018_
rlabel metal1 9384 10438 9384 10438 0 _019_
rlabel metal2 9522 11934 9522 11934 0 _020_
rlabel metal1 10488 12886 10488 12886 0 _021_
rlabel metal2 11086 9316 11086 9316 0 _022_
rlabel metal1 10856 8058 10856 8058 0 _023_
rlabel metal2 8694 5406 8694 5406 0 _024_
rlabel metal1 10902 7174 10902 7174 0 _025_
rlabel metal1 10534 5338 10534 5338 0 _026_
rlabel metal1 10856 2618 10856 2618 0 _027_
rlabel metal1 11185 3094 11185 3094 0 _028_
rlabel metal2 9062 2822 9062 2822 0 _029_
rlabel metal1 4416 10030 4416 10030 0 _030_
rlabel metal1 5750 9146 5750 9146 0 _031_
rlabel metal2 3450 7004 3450 7004 0 _032_
rlabel metal1 2124 6358 2124 6358 0 _033_
rlabel metal1 1978 6834 1978 6834 0 _034_
rlabel metal1 2484 6086 2484 6086 0 _035_
rlabel metal2 3082 5474 3082 5474 0 _036_
rlabel metal2 3266 4250 3266 4250 0 _037_
rlabel metal1 4922 5338 4922 5338 0 _038_
rlabel metal2 5382 4522 5382 4522 0 _039_
rlabel metal1 5842 2924 5842 2924 0 _040_
rlabel metal1 6578 3060 6578 3060 0 _041_
rlabel metal1 6808 3162 6808 3162 0 _042_
rlabel metal1 5704 4250 5704 4250 0 _043_
rlabel metal1 6578 5236 6578 5236 0 _044_
rlabel metal1 7774 8432 7774 8432 0 _045_
rlabel metal1 7590 8500 7590 8500 0 _046_
rlabel metal1 8924 8058 8924 8058 0 _047_
rlabel metal2 8602 10234 8602 10234 0 _048_
rlabel metal1 10718 8602 10718 8602 0 _049_
rlabel metal2 10074 9384 10074 9384 0 _050_
rlabel metal1 10948 12818 10948 12818 0 _051_
rlabel metal1 9890 12308 9890 12308 0 _052_
rlabel metal1 12052 10778 12052 10778 0 _053_
rlabel metal1 9568 7854 9568 7854 0 _054_
rlabel metal1 9430 7888 9430 7888 0 _055_
rlabel metal2 9798 5508 9798 5508 0 _056_
rlabel metal1 10580 5746 10580 5746 0 _057_
rlabel metal1 11170 4454 11170 4454 0 _058_
rlabel metal1 9623 4046 9623 4046 0 _059_
rlabel metal1 10764 4454 10764 4454 0 _060_
rlabel metal1 8970 2482 8970 2482 0 _061_
rlabel metal1 5750 11764 5750 11764 0 _062_
rlabel metal2 5934 11900 5934 11900 0 _063_
rlabel metal2 1978 10540 1978 10540 0 _064_
rlabel metal1 4370 11288 4370 11288 0 _065_
rlabel metal2 4186 9741 4186 9741 0 clk
rlabel metal1 6946 9622 6946 9622 0 clknet_0_clk
rlabel metal1 1932 3570 1932 3570 0 clknet_2_0__leaf_clk
rlabel metal1 9614 6324 9614 6324 0 clknet_2_1__leaf_clk
rlabel metal1 1472 9486 1472 9486 0 clknet_2_2__leaf_clk
rlabel metal2 7038 7616 7038 7616 0 clknet_2_3__leaf_clk
rlabel metal3 751 5508 751 5508 0 current_pc[10]
rlabel metal3 751 6188 751 6188 0 current_pc[11]
rlabel metal2 3266 1520 3266 1520 0 current_pc[12]
rlabel metal2 3910 1520 3910 1520 0 current_pc[13]
rlabel metal2 5842 1520 5842 1520 0 current_pc[14]
rlabel metal2 6486 959 6486 959 0 current_pc[15]
rlabel metal2 7774 1520 7774 1520 0 current_pc[16]
rlabel metal2 7130 1520 7130 1520 0 current_pc[17]
rlabel metal2 11454 7633 11454 7633 0 current_pc[18]
rlabel metal1 11684 8330 11684 8330 0 current_pc[19]
rlabel metal1 11960 8602 11960 8602 0 current_pc[20]
rlabel metal1 11868 11526 11868 11526 0 current_pc[21]
rlabel metal1 10856 12614 10856 12614 0 current_pc[22]
rlabel metal1 11914 12614 11914 12614 0 current_pc[23]
rlabel metal1 11822 10234 11822 10234 0 current_pc[24]
rlabel metal1 11868 8058 11868 8058 0 current_pc[25]
rlabel metal1 11868 4794 11868 4794 0 current_pc[26]
rlabel metal1 11822 7174 11822 7174 0 current_pc[27]
rlabel metal1 11776 4726 11776 4726 0 current_pc[28]
rlabel metal2 11822 4063 11822 4063 0 current_pc[29]
rlabel metal1 4600 12954 4600 12954 0 current_pc[2]
rlabel metal2 11822 3417 11822 3417 0 current_pc[30]
rlabel metal2 9062 1520 9062 1520 0 current_pc[31]
rlabel metal2 5014 13923 5014 13923 0 current_pc[3]
rlabel metal2 6762 13923 6762 13923 0 current_pc[4]
rlabel metal2 6118 13923 6118 13923 0 current_pc[5]
rlabel metal3 751 9588 751 9588 0 current_pc[6]
rlabel metal3 751 8908 751 8908 0 current_pc[7]
rlabel metal3 751 8228 751 8228 0 current_pc[8]
rlabel metal3 751 7548 751 7548 0 current_pc[9]
rlabel metal1 11500 3162 11500 3162 0 net1
rlabel metal1 8740 7514 8740 7514 0 net10
rlabel metal1 11316 9894 11316 9894 0 net11
rlabel metal1 8740 9146 8740 9146 0 net12
rlabel metal2 10994 10914 10994 10914 0 net13
rlabel metal2 11178 11220 11178 11220 0 net14
rlabel metal1 11868 12818 11868 12818 0 net15
rlabel metal1 11408 10778 11408 10778 0 net16
rlabel metal1 11040 8534 11040 8534 0 net17
rlabel metal1 9614 5338 9614 5338 0 net18
rlabel metal1 11730 5032 11730 5032 0 net19
rlabel metal1 1702 5712 1702 5712 0 net2
rlabel metal1 11362 5746 11362 5746 0 net20
rlabel metal1 10488 4114 10488 4114 0 net21
rlabel metal1 4738 12784 4738 12784 0 net22
rlabel metal2 10442 4148 10442 4148 0 net23
rlabel metal1 10074 2414 10074 2414 0 net24
rlabel metal1 5060 12818 5060 12818 0 net25
rlabel metal1 6624 12818 6624 12818 0 net26
rlabel metal1 5980 12818 5980 12818 0 net27
rlabel metal2 2714 10370 2714 10370 0 net28
rlabel metal1 2208 8602 2208 8602 0 net29
rlabel metal1 1932 6086 1932 6086 0 net3
rlabel metal2 2622 8194 2622 8194 0 net30
rlabel metal2 2714 7616 2714 7616 0 net31
rlabel metal1 4554 2380 4554 2380 0 net32
rlabel metal1 11132 2414 11132 2414 0 net33
rlabel metal1 3726 10030 3726 10030 0 net34
rlabel metal1 9890 12818 9890 12818 0 net35
rlabel metal1 11960 2618 11960 2618 0 net36
rlabel metal1 10258 12682 10258 12682 0 net37
rlabel metal1 8602 2380 8602 2380 0 net38
rlabel metal1 10626 5678 10626 5678 0 net39
rlabel metal1 3542 2414 3542 2414 0 net4
rlabel metal1 9338 3502 9338 3502 0 net40
rlabel metal1 4554 12206 4554 12206 0 net41
rlabel metal1 2944 4114 2944 4114 0 net42
rlabel metal2 2806 3468 2806 3468 0 net43
rlabel metal1 6118 3026 6118 3026 0 net44
rlabel metal2 7406 4454 7406 4454 0 net45
rlabel metal2 3266 8636 3266 8636 0 net46
rlabel metal1 11040 12274 11040 12274 0 net47
rlabel metal1 2254 10030 2254 10030 0 net48
rlabel metal1 5612 12818 5612 12818 0 net49
rlabel metal1 4278 2448 4278 2448 0 net5
rlabel metal1 2208 5202 2208 5202 0 net50
rlabel metal2 9798 9826 9798 9826 0 net51
rlabel metal1 7038 5236 7038 5236 0 net52
rlabel metal1 5290 3060 5290 3060 0 net53
rlabel metal1 11454 9554 11454 9554 0 net54
rlabel metal1 9338 11152 9338 11152 0 net55
rlabel metal2 8878 6596 8878 6596 0 net56
rlabel metal1 7912 6766 7912 6766 0 net57
rlabel metal1 8326 8466 8326 8466 0 net58
rlabel metal2 11362 12206 11362 12206 0 net59
rlabel metal1 6210 2448 6210 2448 0 net6
rlabel metal1 9890 4182 9890 4182 0 net60
rlabel metal1 11500 5610 11500 5610 0 net61
rlabel metal2 9154 8330 9154 8330 0 net62
rlabel metal1 6808 2414 6808 2414 0 net7
rlabel metal1 8142 2482 8142 2482 0 net8
rlabel metal1 7406 2414 7406 2414 0 net9
rlabel metal1 11868 3026 11868 3026 0 reset
<< properties >>
string FIXED_BBOX 0 0 120000 120000
<< end >>
